(*use_dsp = "yes"*)
module tdot (
    input wire clock,
    input wire reset,
    input wire [7:0] a0,
    input wire [7:0] c0,
    input wire [7:0] e0,
    input wire [7:0] g0,
    input wire [7:0] i0,
    input wire [7:0] a1,
    input wire [7:0] c1,
    input wire [7:0] e1,
    input wire [7:0] g1,
    input wire [7:0] i1,
    input wire [7:0] a2,
    input wire [7:0] c2,
    input wire [7:0] e2,
    input wire [7:0] g2,
    input wire [7:0] i2,
    input wire [7:0] a3,
    input wire [7:0] c3,
    input wire [7:0] e3,
    input wire [7:0] g3,
    input wire [7:0] i3,
    input wire [7:0] a4,
    input wire [7:0] c4,
    input wire [7:0] e4,
    input wire [7:0] g4,
    input wire [7:0] i4,
    input wire [7:0] a5,
    input wire [7:0] c5,
    input wire [7:0] e5,
    input wire [7:0] g5,
    input wire [7:0] i5,
    input wire [7:0] a6,
    input wire [7:0] c6,
    input wire [7:0] e6,
    input wire [7:0] g6,
    input wire [7:0] i6,
    input wire [7:0] a7,
    input wire [7:0] c7,
    input wire [7:0] e7,
    input wire [7:0] g7,
    input wire [7:0] i7,
    input wire [7:0] a8,
    input wire [7:0] c8,
    input wire [7:0] e8,
    input wire [7:0] g8,
    input wire [7:0] i8,
    input wire [7:0] b0,
    input wire [7:0] d0,
    input wire [7:0] f0,
    input wire [7:0] h0,
    input wire [7:0] j0,
    input wire [7:0] b1,
    input wire [7:0] d1,
    input wire [7:0] f1,
    input wire [7:0] h1,
    input wire [7:0] j1,
    input wire [7:0] b2,
    input wire [7:0] d2,
    input wire [7:0] f2,
    input wire [7:0] h2,
    input wire [7:0] j2,
    input wire [7:0] b3,
    input wire [7:0] d3,
    input wire [7:0] f3,
    input wire [7:0] h3,
    input wire [7:0] j3,
    input wire [7:0] b4,
    input wire [7:0] d4,
    input wire [7:0] f4,
    input wire [7:0] h4,
    input wire [7:0] j4,
    input wire [7:0] b5,
    input wire [7:0] d5,
    input wire [7:0] f5,
    input wire [7:0] h5,
    input wire [7:0] j5,
    input wire [7:0] b6,
    input wire [7:0] d6,
    input wire [7:0] f6,
    input wire [7:0] h6,
    input wire [7:0] j6,
    input wire [7:0] b7,
    input wire [7:0] d7,
    input wire [7:0] f7,
    input wire [7:0] h7,
    input wire [7:0] j7,
    input wire [7:0] b8,
    input wire [7:0] d8,
    input wire [7:0] f8,
    input wire [7:0] h8,
    input wire [7:0] j8,
    input wire [7:0] m,
    input wire [7:0] n,
    input wire [7:0] o,
    input wire [7:0] p,
    input wire [7:0] q,
    input wire en,
    output reg [7:0] v,
    output reg [7:0] w,
    output reg [7:0] x,
    output reg [7:0] y,
    output reg [7:0] z
);
    reg [7:0] t0;
    reg [7:0] t1;
    wire [7:0] t2;
    reg [7:0] t3;
    wire [7:0] t4;
    reg [7:0] t5;
    reg [7:0] t6;
    reg [7:0] t7;
    wire [7:0] t8;
    reg [7:0] t9;
    wire [7:0] t10;
    reg [7:0] t11;
    reg [7:0] t12;
    reg [7:0] t13;
    wire [7:0] t14;
    reg [7:0] t15;
    wire [7:0] t16;
    reg [7:0] t17;
    reg [7:0] t18;
    reg [7:0] t19;
    wire [7:0] t20;
    reg [7:0] t21;
    wire [7:0] t22;
    reg [7:0] t23;
    reg [7:0] t24;
    reg [7:0] t25;
    wire [7:0] t26;
    reg [7:0] t27;
    wire [7:0] t28;
    reg [7:0] t29;
    reg [7:0] t30;
    reg [7:0] t31;
    wire [7:0] t32;
    reg [7:0] t33;
    wire [7:0] t34;
    reg [7:0] t35;
    reg [7:0] t36;
    reg [7:0] t37;
    wire [7:0] t38;
    reg [7:0] t39;
    wire [7:0] t40;
    reg [7:0] t41;
    reg [7:0] t42;
    reg [7:0] t43;
    wire [7:0] t44;
    reg [7:0] t45;
    wire [7:0] t46;
    reg [7:0] t47;
    reg [7:0] t48;
    reg [7:0] t49;
    wire [7:0] t50;
    reg [7:0] t51;
    wire [7:0] t52;
    reg [7:0] t54;
    reg [7:0] t55;
    wire [7:0] t56;
    reg [7:0] t57;
    wire [7:0] t58;
    reg [7:0] t59;
    reg [7:0] t60;
    reg [7:0] t61;
    wire [7:0] t62;
    reg [7:0] t63;
    wire [7:0] t64;
    reg [7:0] t65;
    reg [7:0] t66;
    reg [7:0] t67;
    wire [7:0] t68;
    reg [7:0] t69;
    wire [7:0] t70;
    reg [7:0] t71;
    reg [7:0] t72;
    reg [7:0] t73;
    wire [7:0] t74;
    reg [7:0] t75;
    wire [7:0] t76;
    reg [7:0] t77;
    reg [7:0] t78;
    reg [7:0] t79;
    wire [7:0] t80;
    reg [7:0] t81;
    wire [7:0] t82;
    reg [7:0] t83;
    reg [7:0] t84;
    reg [7:0] t85;
    wire [7:0] t86;
    reg [7:0] t87;
    wire [7:0] t88;
    reg [7:0] t89;
    reg [7:0] t90;
    reg [7:0] t91;
    wire [7:0] t92;
    reg [7:0] t93;
    wire [7:0] t94;
    reg [7:0] t95;
    reg [7:0] t96;
    reg [7:0] t97;
    wire [7:0] t98;
    reg [7:0] t99;
    wire [7:0] t100;
    reg [7:0] t101;
    reg [7:0] t102;
    reg [7:0] t103;
    wire [7:0] t104;
    reg [7:0] t105;
    wire [7:0] t106;
    reg [7:0] t108;
    reg [7:0] t109;
    wire [7:0] t110;
    reg [7:0] t111;
    wire [7:0] t112;
    reg [7:0] t113;
    reg [7:0] t114;
    reg [7:0] t115;
    wire [7:0] t116;
    reg [7:0] t117;
    wire [7:0] t118;
    reg [7:0] t119;
    reg [7:0] t120;
    reg [7:0] t121;
    wire [7:0] t122;
    reg [7:0] t123;
    wire [7:0] t124;
    reg [7:0] t125;
    reg [7:0] t126;
    reg [7:0] t127;
    wire [7:0] t128;
    reg [7:0] t129;
    wire [7:0] t130;
    reg [7:0] t131;
    reg [7:0] t132;
    reg [7:0] t133;
    wire [7:0] t134;
    reg [7:0] t135;
    wire [7:0] t136;
    reg [7:0] t137;
    reg [7:0] t138;
    reg [7:0] t139;
    wire [7:0] t140;
    reg [7:0] t141;
    wire [7:0] t142;
    reg [7:0] t143;
    reg [7:0] t144;
    reg [7:0] t145;
    wire [7:0] t146;
    reg [7:0] t147;
    wire [7:0] t148;
    reg [7:0] t149;
    reg [7:0] t150;
    reg [7:0] t151;
    wire [7:0] t152;
    reg [7:0] t153;
    wire [7:0] t154;
    reg [7:0] t155;
    reg [7:0] t156;
    reg [7:0] t157;
    wire [7:0] t158;
    reg [7:0] t159;
    wire [7:0] t160;
    reg [7:0] t162;
    reg [7:0] t163;
    wire [7:0] t164;
    reg [7:0] t165;
    wire [7:0] t166;
    reg [7:0] t167;
    reg [7:0] t168;
    reg [7:0] t169;
    wire [7:0] t170;
    reg [7:0] t171;
    wire [7:0] t172;
    reg [7:0] t173;
    reg [7:0] t174;
    reg [7:0] t175;
    wire [7:0] t176;
    reg [7:0] t177;
    wire [7:0] t178;
    reg [7:0] t179;
    reg [7:0] t180;
    reg [7:0] t181;
    wire [7:0] t182;
    reg [7:0] t183;
    wire [7:0] t184;
    reg [7:0] t185;
    reg [7:0] t186;
    reg [7:0] t187;
    wire [7:0] t188;
    reg [7:0] t189;
    wire [7:0] t190;
    reg [7:0] t191;
    reg [7:0] t192;
    reg [7:0] t193;
    wire [7:0] t194;
    reg [7:0] t195;
    wire [7:0] t196;
    reg [7:0] t197;
    reg [7:0] t198;
    reg [7:0] t199;
    wire [7:0] t200;
    reg [7:0] t201;
    wire [7:0] t202;
    reg [7:0] t203;
    reg [7:0] t204;
    reg [7:0] t205;
    wire [7:0] t206;
    reg [7:0] t207;
    wire [7:0] t208;
    reg [7:0] t209;
    reg [7:0] t210;
    reg [7:0] t211;
    wire [7:0] t212;
    reg [7:0] t213;
    wire [7:0] t214;
    reg [7:0] t216;
    reg [7:0] t217;
    wire [7:0] t218;
    reg [7:0] t219;
    wire [7:0] t220;
    reg [7:0] t221;
    reg [7:0] t222;
    reg [7:0] t223;
    wire [7:0] t224;
    reg [7:0] t225;
    wire [7:0] t226;
    reg [7:0] t227;
    reg [7:0] t228;
    reg [7:0] t229;
    wire [7:0] t230;
    reg [7:0] t231;
    wire [7:0] t232;
    reg [7:0] t233;
    reg [7:0] t234;
    reg [7:0] t235;
    wire [7:0] t236;
    reg [7:0] t237;
    wire [7:0] t238;
    reg [7:0] t239;
    reg [7:0] t240;
    reg [7:0] t241;
    wire [7:0] t242;
    reg [7:0] t243;
    wire [7:0] t244;
    reg [7:0] t245;
    reg [7:0] t246;
    reg [7:0] t247;
    wire [7:0] t248;
    reg [7:0] t249;
    wire [7:0] t250;
    reg [7:0] t251;
    reg [7:0] t252;
    reg [7:0] t253;
    wire [7:0] t254;
    reg [7:0] t255;
    wire [7:0] t256;
    reg [7:0] t257;
    reg [7:0] t258;
    reg [7:0] t259;
    wire [7:0] t260;
    reg [7:0] t261;
    wire [7:0] t262;
    reg [7:0] t263;
    reg [7:0] t264;
    reg [7:0] t265;
    wire [7:0] t266;
    reg [7:0] t267;
    wire [7:0] t268;
    always @(posedge clock) begin
        if(reset) begin
            t0 <= 0;
        end else if(en) begin
            t0 <= a0;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t1 <= 0;
        end else if(en) begin
            t1 <= b0;
        end
    end
    assign t2 = ($signed(t0) * $signed(t1));
    always @(posedge clock) begin
        if(reset) begin
            t3 <= 0;
        end else if(en) begin
            t3 <= t2;
        end
    end
    assign t4 = ($signed(t3) + $signed(m));
    always @(posedge clock) begin
        if(reset) begin
            t5 <= 0;
        end else if(en) begin
            t5 <= t4;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t6 <= 0;
        end else if(en) begin
            t6 <= a1;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t7 <= 0;
        end else if(en) begin
            t7 <= b1;
        end
    end
    assign t8 = ($signed(t6) * $signed(t7));
    always @(posedge clock) begin
        if(reset) begin
            t9 <= 0;
        end else if(en) begin
            t9 <= t8;
        end
    end
    assign t10 = ($signed(t9) + $signed(t5));
    always @(posedge clock) begin
        if(reset) begin
            t11 <= 0;
        end else if(en) begin
            t11 <= t10;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t12 <= 0;
        end else if(en) begin
            t12 <= a2;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t13 <= 0;
        end else if(en) begin
            t13 <= b2;
        end
    end
    assign t14 = ($signed(t12) * $signed(t13));
    always @(posedge clock) begin
        if(reset) begin
            t15 <= 0;
        end else if(en) begin
            t15 <= t14;
        end
    end
    assign t16 = ($signed(t15) + $signed(t11));
    always @(posedge clock) begin
        if(reset) begin
            t17 <= 0;
        end else if(en) begin
            t17 <= t16;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t18 <= 0;
        end else if(en) begin
            t18 <= a3;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t19 <= 0;
        end else if(en) begin
            t19 <= b3;
        end
    end
    assign t20 = ($signed(t18) * $signed(t19));
    always @(posedge clock) begin
        if(reset) begin
            t21 <= 0;
        end else if(en) begin
            t21 <= t20;
        end
    end
    assign t22 = ($signed(t21) + $signed(t17));
    always @(posedge clock) begin
        if(reset) begin
            t23 <= 0;
        end else if(en) begin
            t23 <= t22;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t24 <= 0;
        end else if(en) begin
            t24 <= a4;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t25 <= 0;
        end else if(en) begin
            t25 <= b4;
        end
    end
    assign t26 = ($signed(t24) * $signed(t25));
    always @(posedge clock) begin
        if(reset) begin
            t27 <= 0;
        end else if(en) begin
            t27 <= t26;
        end
    end
    assign t28 = ($signed(t27) + $signed(t23));
    always @(posedge clock) begin
        if(reset) begin
            t29 <= 0;
        end else if(en) begin
            t29 <= t28;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t30 <= 0;
        end else if(en) begin
            t30 <= a5;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t31 <= 0;
        end else if(en) begin
            t31 <= b5;
        end
    end
    assign t32 = ($signed(t30) * $signed(t31));
    always @(posedge clock) begin
        if(reset) begin
            t33 <= 0;
        end else if(en) begin
            t33 <= t32;
        end
    end
    assign t34 = ($signed(t33) + $signed(t29));
    always @(posedge clock) begin
        if(reset) begin
            t35 <= 0;
        end else if(en) begin
            t35 <= t34;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t36 <= 0;
        end else if(en) begin
            t36 <= a6;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t37 <= 0;
        end else if(en) begin
            t37 <= b6;
        end
    end
    assign t38 = ($signed(t36) * $signed(t37));
    always @(posedge clock) begin
        if(reset) begin
            t39 <= 0;
        end else if(en) begin
            t39 <= t38;
        end
    end
    assign t40 = ($signed(t39) + $signed(t35));
    always @(posedge clock) begin
        if(reset) begin
            t41 <= 0;
        end else if(en) begin
            t41 <= t40;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t42 <= 0;
        end else if(en) begin
            t42 <= a7;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t43 <= 0;
        end else if(en) begin
            t43 <= b7;
        end
    end
    assign t44 = ($signed(t42) * $signed(t43));
    always @(posedge clock) begin
        if(reset) begin
            t45 <= 0;
        end else if(en) begin
            t45 <= t44;
        end
    end
    assign t46 = ($signed(t45) + $signed(t41));
    always @(posedge clock) begin
        if(reset) begin
            t47 <= 0;
        end else if(en) begin
            t47 <= t46;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t48 <= 0;
        end else if(en) begin
            t48 <= a8;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t49 <= 0;
        end else if(en) begin
            t49 <= b8;
        end
    end
    assign t50 = ($signed(t48) * $signed(t49));
    always @(posedge clock) begin
        if(reset) begin
            t51 <= 0;
        end else if(en) begin
            t51 <= t50;
        end
    end
    assign t52 = ($signed(t51) + $signed(t47));
    always @(posedge clock) begin
        if(reset) begin
            v <= 0;
        end else if(en) begin
            v <= t52;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t54 <= 0;
        end else if(en) begin
            t54 <= c0;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t55 <= 0;
        end else if(en) begin
            t55 <= d0;
        end
    end
    assign t56 = ($signed(t54) * $signed(t55));
    always @(posedge clock) begin
        if(reset) begin
            t57 <= 0;
        end else if(en) begin
            t57 <= t56;
        end
    end
    assign t58 = ($signed(t57) + $signed(n));
    always @(posedge clock) begin
        if(reset) begin
            t59 <= 0;
        end else if(en) begin
            t59 <= t58;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t60 <= 0;
        end else if(en) begin
            t60 <= c1;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t61 <= 0;
        end else if(en) begin
            t61 <= d1;
        end
    end
    assign t62 = ($signed(t60) * $signed(t61));
    always @(posedge clock) begin
        if(reset) begin
            t63 <= 0;
        end else if(en) begin
            t63 <= t62;
        end
    end
    assign t64 = ($signed(t63) + $signed(t59));
    always @(posedge clock) begin
        if(reset) begin
            t65 <= 0;
        end else if(en) begin
            t65 <= t64;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t66 <= 0;
        end else if(en) begin
            t66 <= c2;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t67 <= 0;
        end else if(en) begin
            t67 <= d2;
        end
    end
    assign t68 = ($signed(t66) * $signed(t67));
    always @(posedge clock) begin
        if(reset) begin
            t69 <= 0;
        end else if(en) begin
            t69 <= t68;
        end
    end
    assign t70 = ($signed(t69) + $signed(t65));
    always @(posedge clock) begin
        if(reset) begin
            t71 <= 0;
        end else if(en) begin
            t71 <= t70;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t72 <= 0;
        end else if(en) begin
            t72 <= c3;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t73 <= 0;
        end else if(en) begin
            t73 <= d3;
        end
    end
    assign t74 = ($signed(t72) * $signed(t73));
    always @(posedge clock) begin
        if(reset) begin
            t75 <= 0;
        end else if(en) begin
            t75 <= t74;
        end
    end
    assign t76 = ($signed(t75) + $signed(t71));
    always @(posedge clock) begin
        if(reset) begin
            t77 <= 0;
        end else if(en) begin
            t77 <= t76;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t78 <= 0;
        end else if(en) begin
            t78 <= c4;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t79 <= 0;
        end else if(en) begin
            t79 <= d4;
        end
    end
    assign t80 = ($signed(t78) * $signed(t79));
    always @(posedge clock) begin
        if(reset) begin
            t81 <= 0;
        end else if(en) begin
            t81 <= t80;
        end
    end
    assign t82 = ($signed(t81) + $signed(t77));
    always @(posedge clock) begin
        if(reset) begin
            t83 <= 0;
        end else if(en) begin
            t83 <= t82;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t84 <= 0;
        end else if(en) begin
            t84 <= c5;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t85 <= 0;
        end else if(en) begin
            t85 <= d5;
        end
    end
    assign t86 = ($signed(t84) * $signed(t85));
    always @(posedge clock) begin
        if(reset) begin
            t87 <= 0;
        end else if(en) begin
            t87 <= t86;
        end
    end
    assign t88 = ($signed(t87) + $signed(t83));
    always @(posedge clock) begin
        if(reset) begin
            t89 <= 0;
        end else if(en) begin
            t89 <= t88;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t90 <= 0;
        end else if(en) begin
            t90 <= c6;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t91 <= 0;
        end else if(en) begin
            t91 <= d6;
        end
    end
    assign t92 = ($signed(t90) * $signed(t91));
    always @(posedge clock) begin
        if(reset) begin
            t93 <= 0;
        end else if(en) begin
            t93 <= t92;
        end
    end
    assign t94 = ($signed(t93) + $signed(t89));
    always @(posedge clock) begin
        if(reset) begin
            t95 <= 0;
        end else if(en) begin
            t95 <= t94;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t96 <= 0;
        end else if(en) begin
            t96 <= c7;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t97 <= 0;
        end else if(en) begin
            t97 <= d7;
        end
    end
    assign t98 = ($signed(t96) * $signed(t97));
    always @(posedge clock) begin
        if(reset) begin
            t99 <= 0;
        end else if(en) begin
            t99 <= t98;
        end
    end
    assign t100 = ($signed(t99) + $signed(t95));
    always @(posedge clock) begin
        if(reset) begin
            t101 <= 0;
        end else if(en) begin
            t101 <= t100;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t102 <= 0;
        end else if(en) begin
            t102 <= c8;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t103 <= 0;
        end else if(en) begin
            t103 <= d8;
        end
    end
    assign t104 = ($signed(t102) * $signed(t103));
    always @(posedge clock) begin
        if(reset) begin
            t105 <= 0;
        end else if(en) begin
            t105 <= t104;
        end
    end
    assign t106 = ($signed(t105) + $signed(t101));
    always @(posedge clock) begin
        if(reset) begin
            w <= 0;
        end else if(en) begin
            w <= t106;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t108 <= 0;
        end else if(en) begin
            t108 <= e0;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t109 <= 0;
        end else if(en) begin
            t109 <= f0;
        end
    end
    assign t110 = ($signed(t108) * $signed(t109));
    always @(posedge clock) begin
        if(reset) begin
            t111 <= 0;
        end else if(en) begin
            t111 <= t110;
        end
    end
    assign t112 = ($signed(t111) + $signed(o));
    always @(posedge clock) begin
        if(reset) begin
            t113 <= 0;
        end else if(en) begin
            t113 <= t112;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t114 <= 0;
        end else if(en) begin
            t114 <= e1;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t115 <= 0;
        end else if(en) begin
            t115 <= f1;
        end
    end
    assign t116 = ($signed(t114) * $signed(t115));
    always @(posedge clock) begin
        if(reset) begin
            t117 <= 0;
        end else if(en) begin
            t117 <= t116;
        end
    end
    assign t118 = ($signed(t117) + $signed(t113));
    always @(posedge clock) begin
        if(reset) begin
            t119 <= 0;
        end else if(en) begin
            t119 <= t118;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t120 <= 0;
        end else if(en) begin
            t120 <= e2;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t121 <= 0;
        end else if(en) begin
            t121 <= f2;
        end
    end
    assign t122 = ($signed(t120) * $signed(t121));
    always @(posedge clock) begin
        if(reset) begin
            t123 <= 0;
        end else if(en) begin
            t123 <= t122;
        end
    end
    assign t124 = ($signed(t123) + $signed(t119));
    always @(posedge clock) begin
        if(reset) begin
            t125 <= 0;
        end else if(en) begin
            t125 <= t124;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t126 <= 0;
        end else if(en) begin
            t126 <= e3;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t127 <= 0;
        end else if(en) begin
            t127 <= f3;
        end
    end
    assign t128 = ($signed(t126) * $signed(t127));
    always @(posedge clock) begin
        if(reset) begin
            t129 <= 0;
        end else if(en) begin
            t129 <= t128;
        end
    end
    assign t130 = ($signed(t129) + $signed(t125));
    always @(posedge clock) begin
        if(reset) begin
            t131 <= 0;
        end else if(en) begin
            t131 <= t130;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t132 <= 0;
        end else if(en) begin
            t132 <= e4;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t133 <= 0;
        end else if(en) begin
            t133 <= f4;
        end
    end
    assign t134 = ($signed(t132) * $signed(t133));
    always @(posedge clock) begin
        if(reset) begin
            t135 <= 0;
        end else if(en) begin
            t135 <= t134;
        end
    end
    assign t136 = ($signed(t135) + $signed(t131));
    always @(posedge clock) begin
        if(reset) begin
            t137 <= 0;
        end else if(en) begin
            t137 <= t136;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t138 <= 0;
        end else if(en) begin
            t138 <= e5;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t139 <= 0;
        end else if(en) begin
            t139 <= f5;
        end
    end
    assign t140 = ($signed(t138) * $signed(t139));
    always @(posedge clock) begin
        if(reset) begin
            t141 <= 0;
        end else if(en) begin
            t141 <= t140;
        end
    end
    assign t142 = ($signed(t141) + $signed(t137));
    always @(posedge clock) begin
        if(reset) begin
            t143 <= 0;
        end else if(en) begin
            t143 <= t142;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t144 <= 0;
        end else if(en) begin
            t144 <= e6;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t145 <= 0;
        end else if(en) begin
            t145 <= f6;
        end
    end
    assign t146 = ($signed(t144) * $signed(t145));
    always @(posedge clock) begin
        if(reset) begin
            t147 <= 0;
        end else if(en) begin
            t147 <= t146;
        end
    end
    assign t148 = ($signed(t147) + $signed(t143));
    always @(posedge clock) begin
        if(reset) begin
            t149 <= 0;
        end else if(en) begin
            t149 <= t148;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t150 <= 0;
        end else if(en) begin
            t150 <= e7;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t151 <= 0;
        end else if(en) begin
            t151 <= f7;
        end
    end
    assign t152 = ($signed(t150) * $signed(t151));
    always @(posedge clock) begin
        if(reset) begin
            t153 <= 0;
        end else if(en) begin
            t153 <= t152;
        end
    end
    assign t154 = ($signed(t153) + $signed(t149));
    always @(posedge clock) begin
        if(reset) begin
            t155 <= 0;
        end else if(en) begin
            t155 <= t154;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t156 <= 0;
        end else if(en) begin
            t156 <= e8;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t157 <= 0;
        end else if(en) begin
            t157 <= f8;
        end
    end
    assign t158 = ($signed(t156) * $signed(t157));
    always @(posedge clock) begin
        if(reset) begin
            t159 <= 0;
        end else if(en) begin
            t159 <= t158;
        end
    end
    assign t160 = ($signed(t159) + $signed(t155));
    always @(posedge clock) begin
        if(reset) begin
            x <= 0;
        end else if(en) begin
            x <= t160;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t162 <= 0;
        end else if(en) begin
            t162 <= g0;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t163 <= 0;
        end else if(en) begin
            t163 <= h0;
        end
    end
    assign t164 = ($signed(t162) * $signed(t163));
    always @(posedge clock) begin
        if(reset) begin
            t165 <= 0;
        end else if(en) begin
            t165 <= t164;
        end
    end
    assign t166 = ($signed(t165) + $signed(p));
    always @(posedge clock) begin
        if(reset) begin
            t167 <= 0;
        end else if(en) begin
            t167 <= t166;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t168 <= 0;
        end else if(en) begin
            t168 <= g1;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t169 <= 0;
        end else if(en) begin
            t169 <= h1;
        end
    end
    assign t170 = ($signed(t168) * $signed(t169));
    always @(posedge clock) begin
        if(reset) begin
            t171 <= 0;
        end else if(en) begin
            t171 <= t170;
        end
    end
    assign t172 = ($signed(t171) + $signed(t167));
    always @(posedge clock) begin
        if(reset) begin
            t173 <= 0;
        end else if(en) begin
            t173 <= t172;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t174 <= 0;
        end else if(en) begin
            t174 <= g2;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t175 <= 0;
        end else if(en) begin
            t175 <= h2;
        end
    end
    assign t176 = ($signed(t174) * $signed(t175));
    always @(posedge clock) begin
        if(reset) begin
            t177 <= 0;
        end else if(en) begin
            t177 <= t176;
        end
    end
    assign t178 = ($signed(t177) + $signed(t173));
    always @(posedge clock) begin
        if(reset) begin
            t179 <= 0;
        end else if(en) begin
            t179 <= t178;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t180 <= 0;
        end else if(en) begin
            t180 <= g3;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t181 <= 0;
        end else if(en) begin
            t181 <= h3;
        end
    end
    assign t182 = ($signed(t180) * $signed(t181));
    always @(posedge clock) begin
        if(reset) begin
            t183 <= 0;
        end else if(en) begin
            t183 <= t182;
        end
    end
    assign t184 = ($signed(t183) + $signed(t179));
    always @(posedge clock) begin
        if(reset) begin
            t185 <= 0;
        end else if(en) begin
            t185 <= t184;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t186 <= 0;
        end else if(en) begin
            t186 <= g4;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t187 <= 0;
        end else if(en) begin
            t187 <= h4;
        end
    end
    assign t188 = ($signed(t186) * $signed(t187));
    always @(posedge clock) begin
        if(reset) begin
            t189 <= 0;
        end else if(en) begin
            t189 <= t188;
        end
    end
    assign t190 = ($signed(t189) + $signed(t185));
    always @(posedge clock) begin
        if(reset) begin
            t191 <= 0;
        end else if(en) begin
            t191 <= t190;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t192 <= 0;
        end else if(en) begin
            t192 <= g5;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t193 <= 0;
        end else if(en) begin
            t193 <= h5;
        end
    end
    assign t194 = ($signed(t192) * $signed(t193));
    always @(posedge clock) begin
        if(reset) begin
            t195 <= 0;
        end else if(en) begin
            t195 <= t194;
        end
    end
    assign t196 = ($signed(t195) + $signed(t191));
    always @(posedge clock) begin
        if(reset) begin
            t197 <= 0;
        end else if(en) begin
            t197 <= t196;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t198 <= 0;
        end else if(en) begin
            t198 <= g6;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t199 <= 0;
        end else if(en) begin
            t199 <= h6;
        end
    end
    assign t200 = ($signed(t198) * $signed(t199));
    always @(posedge clock) begin
        if(reset) begin
            t201 <= 0;
        end else if(en) begin
            t201 <= t200;
        end
    end
    assign t202 = ($signed(t201) + $signed(t197));
    always @(posedge clock) begin
        if(reset) begin
            t203 <= 0;
        end else if(en) begin
            t203 <= t202;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t204 <= 0;
        end else if(en) begin
            t204 <= g7;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t205 <= 0;
        end else if(en) begin
            t205 <= h7;
        end
    end
    assign t206 = ($signed(t204) * $signed(t205));
    always @(posedge clock) begin
        if(reset) begin
            t207 <= 0;
        end else if(en) begin
            t207 <= t206;
        end
    end
    assign t208 = ($signed(t207) + $signed(t203));
    always @(posedge clock) begin
        if(reset) begin
            t209 <= 0;
        end else if(en) begin
            t209 <= t208;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t210 <= 0;
        end else if(en) begin
            t210 <= g8;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t211 <= 0;
        end else if(en) begin
            t211 <= h8;
        end
    end
    assign t212 = ($signed(t210) * $signed(t211));
    always @(posedge clock) begin
        if(reset) begin
            t213 <= 0;
        end else if(en) begin
            t213 <= t212;
        end
    end
    assign t214 = ($signed(t213) + $signed(t209));
    always @(posedge clock) begin
        if(reset) begin
            y <= 0;
        end else if(en) begin
            y <= t214;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t216 <= 0;
        end else if(en) begin
            t216 <= i0;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t217 <= 0;
        end else if(en) begin
            t217 <= j0;
        end
    end
    assign t218 = ($signed(t216) * $signed(t217));
    always @(posedge clock) begin
        if(reset) begin
            t219 <= 0;
        end else if(en) begin
            t219 <= t218;
        end
    end
    assign t220 = ($signed(t219) + $signed(q));
    always @(posedge clock) begin
        if(reset) begin
            t221 <= 0;
        end else if(en) begin
            t221 <= t220;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t222 <= 0;
        end else if(en) begin
            t222 <= i1;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t223 <= 0;
        end else if(en) begin
            t223 <= j1;
        end
    end
    assign t224 = ($signed(t222) * $signed(t223));
    always @(posedge clock) begin
        if(reset) begin
            t225 <= 0;
        end else if(en) begin
            t225 <= t224;
        end
    end
    assign t226 = ($signed(t225) + $signed(t221));
    always @(posedge clock) begin
        if(reset) begin
            t227 <= 0;
        end else if(en) begin
            t227 <= t226;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t228 <= 0;
        end else if(en) begin
            t228 <= i2;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t229 <= 0;
        end else if(en) begin
            t229 <= j2;
        end
    end
    assign t230 = ($signed(t228) * $signed(t229));
    always @(posedge clock) begin
        if(reset) begin
            t231 <= 0;
        end else if(en) begin
            t231 <= t230;
        end
    end
    assign t232 = ($signed(t231) + $signed(t227));
    always @(posedge clock) begin
        if(reset) begin
            t233 <= 0;
        end else if(en) begin
            t233 <= t232;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t234 <= 0;
        end else if(en) begin
            t234 <= i3;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t235 <= 0;
        end else if(en) begin
            t235 <= j3;
        end
    end
    assign t236 = ($signed(t234) * $signed(t235));
    always @(posedge clock) begin
        if(reset) begin
            t237 <= 0;
        end else if(en) begin
            t237 <= t236;
        end
    end
    assign t238 = ($signed(t237) + $signed(t233));
    always @(posedge clock) begin
        if(reset) begin
            t239 <= 0;
        end else if(en) begin
            t239 <= t238;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t240 <= 0;
        end else if(en) begin
            t240 <= i4;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t241 <= 0;
        end else if(en) begin
            t241 <= j4;
        end
    end
    assign t242 = ($signed(t240) * $signed(t241));
    always @(posedge clock) begin
        if(reset) begin
            t243 <= 0;
        end else if(en) begin
            t243 <= t242;
        end
    end
    assign t244 = ($signed(t243) + $signed(t239));
    always @(posedge clock) begin
        if(reset) begin
            t245 <= 0;
        end else if(en) begin
            t245 <= t244;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t246 <= 0;
        end else if(en) begin
            t246 <= i5;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t247 <= 0;
        end else if(en) begin
            t247 <= j5;
        end
    end
    assign t248 = ($signed(t246) * $signed(t247));
    always @(posedge clock) begin
        if(reset) begin
            t249 <= 0;
        end else if(en) begin
            t249 <= t248;
        end
    end
    assign t250 = ($signed(t249) + $signed(t245));
    always @(posedge clock) begin
        if(reset) begin
            t251 <= 0;
        end else if(en) begin
            t251 <= t250;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t252 <= 0;
        end else if(en) begin
            t252 <= i6;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t253 <= 0;
        end else if(en) begin
            t253 <= j6;
        end
    end
    assign t254 = ($signed(t252) * $signed(t253));
    always @(posedge clock) begin
        if(reset) begin
            t255 <= 0;
        end else if(en) begin
            t255 <= t254;
        end
    end
    assign t256 = ($signed(t255) + $signed(t251));
    always @(posedge clock) begin
        if(reset) begin
            t257 <= 0;
        end else if(en) begin
            t257 <= t256;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t258 <= 0;
        end else if(en) begin
            t258 <= i7;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t259 <= 0;
        end else if(en) begin
            t259 <= j7;
        end
    end
    assign t260 = ($signed(t258) * $signed(t259));
    always @(posedge clock) begin
        if(reset) begin
            t261 <= 0;
        end else if(en) begin
            t261 <= t260;
        end
    end
    assign t262 = ($signed(t261) + $signed(t257));
    always @(posedge clock) begin
        if(reset) begin
            t263 <= 0;
        end else if(en) begin
            t263 <= t262;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t264 <= 0;
        end else if(en) begin
            t264 <= i8;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t265 <= 0;
        end else if(en) begin
            t265 <= j8;
        end
    end
    assign t266 = ($signed(t264) * $signed(t265));
    always @(posedge clock) begin
        if(reset) begin
            t267 <= 0;
        end else if(en) begin
            t267 <= t266;
        end
    end
    assign t268 = ($signed(t267) + $signed(t263));
    always @(posedge clock) begin
        if(reset) begin
            z <= 0;
        end else if(en) begin
            z <= t268;
        end
    end
endmodule
