(*use_dsp = "yes"*)
module tdot (
    input wire clock,
    input wire reset,
    input wire [7:0] a0,
    input wire [7:0] c0,
    input wire [7:0] e0,
    input wire [7:0] g0,
    input wire [7:0] i0,
    input wire [7:0] a1,
    input wire [7:0] c1,
    input wire [7:0] e1,
    input wire [7:0] g1,
    input wire [7:0] i1,
    input wire [7:0] a2,
    input wire [7:0] c2,
    input wire [7:0] e2,
    input wire [7:0] g2,
    input wire [7:0] i2,
    input wire [7:0] a3,
    input wire [7:0] c3,
    input wire [7:0] e3,
    input wire [7:0] g3,
    input wire [7:0] i3,
    input wire [7:0] a4,
    input wire [7:0] c4,
    input wire [7:0] e4,
    input wire [7:0] g4,
    input wire [7:0] i4,
    input wire [7:0] a5,
    input wire [7:0] c5,
    input wire [7:0] e5,
    input wire [7:0] g5,
    input wire [7:0] i5,
    input wire [7:0] a6,
    input wire [7:0] c6,
    input wire [7:0] e6,
    input wire [7:0] g6,
    input wire [7:0] i6,
    input wire [7:0] a7,
    input wire [7:0] c7,
    input wire [7:0] e7,
    input wire [7:0] g7,
    input wire [7:0] i7,
    input wire [7:0] a8,
    input wire [7:0] c8,
    input wire [7:0] e8,
    input wire [7:0] g8,
    input wire [7:0] i8,
    input wire [7:0] a9,
    input wire [7:0] c9,
    input wire [7:0] e9,
    input wire [7:0] g9,
    input wire [7:0] i9,
    input wire [7:0] a10,
    input wire [7:0] c10,
    input wire [7:0] e10,
    input wire [7:0] g10,
    input wire [7:0] i10,
    input wire [7:0] a11,
    input wire [7:0] c11,
    input wire [7:0] e11,
    input wire [7:0] g11,
    input wire [7:0] i11,
    input wire [7:0] a12,
    input wire [7:0] c12,
    input wire [7:0] e12,
    input wire [7:0] g12,
    input wire [7:0] i12,
    input wire [7:0] a13,
    input wire [7:0] c13,
    input wire [7:0] e13,
    input wire [7:0] g13,
    input wire [7:0] i13,
    input wire [7:0] a14,
    input wire [7:0] c14,
    input wire [7:0] e14,
    input wire [7:0] g14,
    input wire [7:0] i14,
    input wire [7:0] a15,
    input wire [7:0] c15,
    input wire [7:0] e15,
    input wire [7:0] g15,
    input wire [7:0] i15,
    input wire [7:0] a16,
    input wire [7:0] c16,
    input wire [7:0] e16,
    input wire [7:0] g16,
    input wire [7:0] i16,
    input wire [7:0] a17,
    input wire [7:0] c17,
    input wire [7:0] e17,
    input wire [7:0] g17,
    input wire [7:0] i17,
    input wire [7:0] b0,
    input wire [7:0] d0,
    input wire [7:0] f0,
    input wire [7:0] h0,
    input wire [7:0] j0,
    input wire [7:0] b1,
    input wire [7:0] d1,
    input wire [7:0] f1,
    input wire [7:0] h1,
    input wire [7:0] j1,
    input wire [7:0] b2,
    input wire [7:0] d2,
    input wire [7:0] f2,
    input wire [7:0] h2,
    input wire [7:0] j2,
    input wire [7:0] b3,
    input wire [7:0] d3,
    input wire [7:0] f3,
    input wire [7:0] h3,
    input wire [7:0] j3,
    input wire [7:0] b4,
    input wire [7:0] d4,
    input wire [7:0] f4,
    input wire [7:0] h4,
    input wire [7:0] j4,
    input wire [7:0] b5,
    input wire [7:0] d5,
    input wire [7:0] f5,
    input wire [7:0] h5,
    input wire [7:0] j5,
    input wire [7:0] b6,
    input wire [7:0] d6,
    input wire [7:0] f6,
    input wire [7:0] h6,
    input wire [7:0] j6,
    input wire [7:0] b7,
    input wire [7:0] d7,
    input wire [7:0] f7,
    input wire [7:0] h7,
    input wire [7:0] j7,
    input wire [7:0] b8,
    input wire [7:0] d8,
    input wire [7:0] f8,
    input wire [7:0] h8,
    input wire [7:0] j8,
    input wire [7:0] b9,
    input wire [7:0] d9,
    input wire [7:0] f9,
    input wire [7:0] h9,
    input wire [7:0] j9,
    input wire [7:0] b10,
    input wire [7:0] d10,
    input wire [7:0] f10,
    input wire [7:0] h10,
    input wire [7:0] j10,
    input wire [7:0] b11,
    input wire [7:0] d11,
    input wire [7:0] f11,
    input wire [7:0] h11,
    input wire [7:0] j11,
    input wire [7:0] b12,
    input wire [7:0] d12,
    input wire [7:0] f12,
    input wire [7:0] h12,
    input wire [7:0] j12,
    input wire [7:0] b13,
    input wire [7:0] d13,
    input wire [7:0] f13,
    input wire [7:0] h13,
    input wire [7:0] j13,
    input wire [7:0] b14,
    input wire [7:0] d14,
    input wire [7:0] f14,
    input wire [7:0] h14,
    input wire [7:0] j14,
    input wire [7:0] b15,
    input wire [7:0] d15,
    input wire [7:0] f15,
    input wire [7:0] h15,
    input wire [7:0] j15,
    input wire [7:0] b16,
    input wire [7:0] d16,
    input wire [7:0] f16,
    input wire [7:0] h16,
    input wire [7:0] j16,
    input wire [7:0] b17,
    input wire [7:0] d17,
    input wire [7:0] f17,
    input wire [7:0] h17,
    input wire [7:0] j17,
    input wire [7:0] m,
    input wire [7:0] n,
    input wire [7:0] o,
    input wire [7:0] p,
    input wire [7:0] q,
    input wire en,
    output reg [7:0] v,
    output reg [7:0] w,
    output reg [7:0] x,
    output reg [7:0] y,
    output reg [7:0] z
);
    reg [7:0] t0;
    reg [7:0] t1;
    wire [7:0] t2;
    reg [7:0] t3;
    wire [7:0] t4;
    reg [7:0] t5;
    reg [7:0] t6;
    reg [7:0] t7;
    wire [7:0] t8;
    reg [7:0] t9;
    wire [7:0] t10;
    reg [7:0] t11;
    reg [7:0] t12;
    reg [7:0] t13;
    wire [7:0] t14;
    reg [7:0] t15;
    wire [7:0] t16;
    reg [7:0] t17;
    reg [7:0] t18;
    reg [7:0] t19;
    wire [7:0] t20;
    reg [7:0] t21;
    wire [7:0] t22;
    reg [7:0] t23;
    reg [7:0] t24;
    reg [7:0] t25;
    wire [7:0] t26;
    reg [7:0] t27;
    wire [7:0] t28;
    reg [7:0] t29;
    reg [7:0] t30;
    reg [7:0] t31;
    wire [7:0] t32;
    reg [7:0] t33;
    wire [7:0] t34;
    reg [7:0] t35;
    reg [7:0] t36;
    reg [7:0] t37;
    wire [7:0] t38;
    reg [7:0] t39;
    wire [7:0] t40;
    reg [7:0] t41;
    reg [7:0] t42;
    reg [7:0] t43;
    wire [7:0] t44;
    reg [7:0] t45;
    wire [7:0] t46;
    reg [7:0] t47;
    reg [7:0] t48;
    reg [7:0] t49;
    wire [7:0] t50;
    reg [7:0] t51;
    wire [7:0] t52;
    reg [7:0] t53;
    reg [7:0] t54;
    reg [7:0] t55;
    wire [7:0] t56;
    reg [7:0] t57;
    wire [7:0] t58;
    reg [7:0] t59;
    reg [7:0] t60;
    reg [7:0] t61;
    wire [7:0] t62;
    reg [7:0] t63;
    wire [7:0] t64;
    reg [7:0] t65;
    reg [7:0] t66;
    reg [7:0] t67;
    wire [7:0] t68;
    reg [7:0] t69;
    wire [7:0] t70;
    reg [7:0] t71;
    reg [7:0] t72;
    reg [7:0] t73;
    wire [7:0] t74;
    reg [7:0] t75;
    wire [7:0] t76;
    reg [7:0] t77;
    reg [7:0] t78;
    reg [7:0] t79;
    wire [7:0] t80;
    reg [7:0] t81;
    wire [7:0] t82;
    reg [7:0] t83;
    reg [7:0] t84;
    reg [7:0] t85;
    wire [7:0] t86;
    reg [7:0] t87;
    wire [7:0] t88;
    reg [7:0] t89;
    reg [7:0] t90;
    reg [7:0] t91;
    wire [7:0] t92;
    reg [7:0] t93;
    wire [7:0] t94;
    reg [7:0] t95;
    reg [7:0] t96;
    reg [7:0] t97;
    wire [7:0] t98;
    reg [7:0] t99;
    wire [7:0] t100;
    reg [7:0] t101;
    reg [7:0] t102;
    reg [7:0] t103;
    wire [7:0] t104;
    reg [7:0] t105;
    wire [7:0] t106;
    reg [7:0] t108;
    reg [7:0] t109;
    wire [7:0] t110;
    reg [7:0] t111;
    wire [7:0] t112;
    reg [7:0] t113;
    reg [7:0] t114;
    reg [7:0] t115;
    wire [7:0] t116;
    reg [7:0] t117;
    wire [7:0] t118;
    reg [7:0] t119;
    reg [7:0] t120;
    reg [7:0] t121;
    wire [7:0] t122;
    reg [7:0] t123;
    wire [7:0] t124;
    reg [7:0] t125;
    reg [7:0] t126;
    reg [7:0] t127;
    wire [7:0] t128;
    reg [7:0] t129;
    wire [7:0] t130;
    reg [7:0] t131;
    reg [7:0] t132;
    reg [7:0] t133;
    wire [7:0] t134;
    reg [7:0] t135;
    wire [7:0] t136;
    reg [7:0] t137;
    reg [7:0] t138;
    reg [7:0] t139;
    wire [7:0] t140;
    reg [7:0] t141;
    wire [7:0] t142;
    reg [7:0] t143;
    reg [7:0] t144;
    reg [7:0] t145;
    wire [7:0] t146;
    reg [7:0] t147;
    wire [7:0] t148;
    reg [7:0] t149;
    reg [7:0] t150;
    reg [7:0] t151;
    wire [7:0] t152;
    reg [7:0] t153;
    wire [7:0] t154;
    reg [7:0] t155;
    reg [7:0] t156;
    reg [7:0] t157;
    wire [7:0] t158;
    reg [7:0] t159;
    wire [7:0] t160;
    reg [7:0] t161;
    reg [7:0] t162;
    reg [7:0] t163;
    wire [7:0] t164;
    reg [7:0] t165;
    wire [7:0] t166;
    reg [7:0] t167;
    reg [7:0] t168;
    reg [7:0] t169;
    wire [7:0] t170;
    reg [7:0] t171;
    wire [7:0] t172;
    reg [7:0] t173;
    reg [7:0] t174;
    reg [7:0] t175;
    wire [7:0] t176;
    reg [7:0] t177;
    wire [7:0] t178;
    reg [7:0] t179;
    reg [7:0] t180;
    reg [7:0] t181;
    wire [7:0] t182;
    reg [7:0] t183;
    wire [7:0] t184;
    reg [7:0] t185;
    reg [7:0] t186;
    reg [7:0] t187;
    wire [7:0] t188;
    reg [7:0] t189;
    wire [7:0] t190;
    reg [7:0] t191;
    reg [7:0] t192;
    reg [7:0] t193;
    wire [7:0] t194;
    reg [7:0] t195;
    wire [7:0] t196;
    reg [7:0] t197;
    reg [7:0] t198;
    reg [7:0] t199;
    wire [7:0] t200;
    reg [7:0] t201;
    wire [7:0] t202;
    reg [7:0] t203;
    reg [7:0] t204;
    reg [7:0] t205;
    wire [7:0] t206;
    reg [7:0] t207;
    wire [7:0] t208;
    reg [7:0] t209;
    reg [7:0] t210;
    reg [7:0] t211;
    wire [7:0] t212;
    reg [7:0] t213;
    wire [7:0] t214;
    reg [7:0] t216;
    reg [7:0] t217;
    wire [7:0] t218;
    reg [7:0] t219;
    wire [7:0] t220;
    reg [7:0] t221;
    reg [7:0] t222;
    reg [7:0] t223;
    wire [7:0] t224;
    reg [7:0] t225;
    wire [7:0] t226;
    reg [7:0] t227;
    reg [7:0] t228;
    reg [7:0] t229;
    wire [7:0] t230;
    reg [7:0] t231;
    wire [7:0] t232;
    reg [7:0] t233;
    reg [7:0] t234;
    reg [7:0] t235;
    wire [7:0] t236;
    reg [7:0] t237;
    wire [7:0] t238;
    reg [7:0] t239;
    reg [7:0] t240;
    reg [7:0] t241;
    wire [7:0] t242;
    reg [7:0] t243;
    wire [7:0] t244;
    reg [7:0] t245;
    reg [7:0] t246;
    reg [7:0] t247;
    wire [7:0] t248;
    reg [7:0] t249;
    wire [7:0] t250;
    reg [7:0] t251;
    reg [7:0] t252;
    reg [7:0] t253;
    wire [7:0] t254;
    reg [7:0] t255;
    wire [7:0] t256;
    reg [7:0] t257;
    reg [7:0] t258;
    reg [7:0] t259;
    wire [7:0] t260;
    reg [7:0] t261;
    wire [7:0] t262;
    reg [7:0] t263;
    reg [7:0] t264;
    reg [7:0] t265;
    wire [7:0] t266;
    reg [7:0] t267;
    wire [7:0] t268;
    reg [7:0] t269;
    reg [7:0] t270;
    reg [7:0] t271;
    wire [7:0] t272;
    reg [7:0] t273;
    wire [7:0] t274;
    reg [7:0] t275;
    reg [7:0] t276;
    reg [7:0] t277;
    wire [7:0] t278;
    reg [7:0] t279;
    wire [7:0] t280;
    reg [7:0] t281;
    reg [7:0] t282;
    reg [7:0] t283;
    wire [7:0] t284;
    reg [7:0] t285;
    wire [7:0] t286;
    reg [7:0] t287;
    reg [7:0] t288;
    reg [7:0] t289;
    wire [7:0] t290;
    reg [7:0] t291;
    wire [7:0] t292;
    reg [7:0] t293;
    reg [7:0] t294;
    reg [7:0] t295;
    wire [7:0] t296;
    reg [7:0] t297;
    wire [7:0] t298;
    reg [7:0] t299;
    reg [7:0] t300;
    reg [7:0] t301;
    wire [7:0] t302;
    reg [7:0] t303;
    wire [7:0] t304;
    reg [7:0] t305;
    reg [7:0] t306;
    reg [7:0] t307;
    wire [7:0] t308;
    reg [7:0] t309;
    wire [7:0] t310;
    reg [7:0] t311;
    reg [7:0] t312;
    reg [7:0] t313;
    wire [7:0] t314;
    reg [7:0] t315;
    wire [7:0] t316;
    reg [7:0] t317;
    reg [7:0] t318;
    reg [7:0] t319;
    wire [7:0] t320;
    reg [7:0] t321;
    wire [7:0] t322;
    reg [7:0] t324;
    reg [7:0] t325;
    wire [7:0] t326;
    reg [7:0] t327;
    wire [7:0] t328;
    reg [7:0] t329;
    reg [7:0] t330;
    reg [7:0] t331;
    wire [7:0] t332;
    reg [7:0] t333;
    wire [7:0] t334;
    reg [7:0] t335;
    reg [7:0] t336;
    reg [7:0] t337;
    wire [7:0] t338;
    reg [7:0] t339;
    wire [7:0] t340;
    reg [7:0] t341;
    reg [7:0] t342;
    reg [7:0] t343;
    wire [7:0] t344;
    reg [7:0] t345;
    wire [7:0] t346;
    reg [7:0] t347;
    reg [7:0] t348;
    reg [7:0] t349;
    wire [7:0] t350;
    reg [7:0] t351;
    wire [7:0] t352;
    reg [7:0] t353;
    reg [7:0] t354;
    reg [7:0] t355;
    wire [7:0] t356;
    reg [7:0] t357;
    wire [7:0] t358;
    reg [7:0] t359;
    reg [7:0] t360;
    reg [7:0] t361;
    wire [7:0] t362;
    reg [7:0] t363;
    wire [7:0] t364;
    reg [7:0] t365;
    reg [7:0] t366;
    reg [7:0] t367;
    wire [7:0] t368;
    reg [7:0] t369;
    wire [7:0] t370;
    reg [7:0] t371;
    reg [7:0] t372;
    reg [7:0] t373;
    wire [7:0] t374;
    reg [7:0] t375;
    wire [7:0] t376;
    reg [7:0] t377;
    reg [7:0] t378;
    reg [7:0] t379;
    wire [7:0] t380;
    reg [7:0] t381;
    wire [7:0] t382;
    reg [7:0] t383;
    reg [7:0] t384;
    reg [7:0] t385;
    wire [7:0] t386;
    reg [7:0] t387;
    wire [7:0] t388;
    reg [7:0] t389;
    reg [7:0] t390;
    reg [7:0] t391;
    wire [7:0] t392;
    reg [7:0] t393;
    wire [7:0] t394;
    reg [7:0] t395;
    reg [7:0] t396;
    reg [7:0] t397;
    wire [7:0] t398;
    reg [7:0] t399;
    wire [7:0] t400;
    reg [7:0] t401;
    reg [7:0] t402;
    reg [7:0] t403;
    wire [7:0] t404;
    reg [7:0] t405;
    wire [7:0] t406;
    reg [7:0] t407;
    reg [7:0] t408;
    reg [7:0] t409;
    wire [7:0] t410;
    reg [7:0] t411;
    wire [7:0] t412;
    reg [7:0] t413;
    reg [7:0] t414;
    reg [7:0] t415;
    wire [7:0] t416;
    reg [7:0] t417;
    wire [7:0] t418;
    reg [7:0] t419;
    reg [7:0] t420;
    reg [7:0] t421;
    wire [7:0] t422;
    reg [7:0] t423;
    wire [7:0] t424;
    reg [7:0] t425;
    reg [7:0] t426;
    reg [7:0] t427;
    wire [7:0] t428;
    reg [7:0] t429;
    wire [7:0] t430;
    reg [7:0] t432;
    reg [7:0] t433;
    wire [7:0] t434;
    reg [7:0] t435;
    wire [7:0] t436;
    reg [7:0] t437;
    reg [7:0] t438;
    reg [7:0] t439;
    wire [7:0] t440;
    reg [7:0] t441;
    wire [7:0] t442;
    reg [7:0] t443;
    reg [7:0] t444;
    reg [7:0] t445;
    wire [7:0] t446;
    reg [7:0] t447;
    wire [7:0] t448;
    reg [7:0] t449;
    reg [7:0] t450;
    reg [7:0] t451;
    wire [7:0] t452;
    reg [7:0] t453;
    wire [7:0] t454;
    reg [7:0] t455;
    reg [7:0] t456;
    reg [7:0] t457;
    wire [7:0] t458;
    reg [7:0] t459;
    wire [7:0] t460;
    reg [7:0] t461;
    reg [7:0] t462;
    reg [7:0] t463;
    wire [7:0] t464;
    reg [7:0] t465;
    wire [7:0] t466;
    reg [7:0] t467;
    reg [7:0] t468;
    reg [7:0] t469;
    wire [7:0] t470;
    reg [7:0] t471;
    wire [7:0] t472;
    reg [7:0] t473;
    reg [7:0] t474;
    reg [7:0] t475;
    wire [7:0] t476;
    reg [7:0] t477;
    wire [7:0] t478;
    reg [7:0] t479;
    reg [7:0] t480;
    reg [7:0] t481;
    wire [7:0] t482;
    reg [7:0] t483;
    wire [7:0] t484;
    reg [7:0] t485;
    reg [7:0] t486;
    reg [7:0] t487;
    wire [7:0] t488;
    reg [7:0] t489;
    wire [7:0] t490;
    reg [7:0] t491;
    reg [7:0] t492;
    reg [7:0] t493;
    wire [7:0] t494;
    reg [7:0] t495;
    wire [7:0] t496;
    reg [7:0] t497;
    reg [7:0] t498;
    reg [7:0] t499;
    wire [7:0] t500;
    reg [7:0] t501;
    wire [7:0] t502;
    reg [7:0] t503;
    reg [7:0] t504;
    reg [7:0] t505;
    wire [7:0] t506;
    reg [7:0] t507;
    wire [7:0] t508;
    reg [7:0] t509;
    reg [7:0] t510;
    reg [7:0] t511;
    wire [7:0] t512;
    reg [7:0] t513;
    wire [7:0] t514;
    reg [7:0] t515;
    reg [7:0] t516;
    reg [7:0] t517;
    wire [7:0] t518;
    reg [7:0] t519;
    wire [7:0] t520;
    reg [7:0] t521;
    reg [7:0] t522;
    reg [7:0] t523;
    wire [7:0] t524;
    reg [7:0] t525;
    wire [7:0] t526;
    reg [7:0] t527;
    reg [7:0] t528;
    reg [7:0] t529;
    wire [7:0] t530;
    reg [7:0] t531;
    wire [7:0] t532;
    reg [7:0] t533;
    reg [7:0] t534;
    reg [7:0] t535;
    wire [7:0] t536;
    reg [7:0] t537;
    wire [7:0] t538;
    always @(posedge clock) begin
        if(reset) begin
            t0 <= 0;
        end else if(en) begin
            t0 <= a0;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t1 <= 0;
        end else if(en) begin
            t1 <= b0;
        end
    end
    assign t2 = ($signed(t0) * $signed(t1));
    always @(posedge clock) begin
        if(reset) begin
            t3 <= 0;
        end else if(en) begin
            t3 <= t2;
        end
    end
    assign t4 = ($signed(t3) + $signed(m));
    always @(posedge clock) begin
        if(reset) begin
            t5 <= 0;
        end else if(en) begin
            t5 <= t4;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t6 <= 0;
        end else if(en) begin
            t6 <= a1;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t7 <= 0;
        end else if(en) begin
            t7 <= b1;
        end
    end
    assign t8 = ($signed(t6) * $signed(t7));
    always @(posedge clock) begin
        if(reset) begin
            t9 <= 0;
        end else if(en) begin
            t9 <= t8;
        end
    end
    assign t10 = ($signed(t9) + $signed(t5));
    always @(posedge clock) begin
        if(reset) begin
            t11 <= 0;
        end else if(en) begin
            t11 <= t10;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t12 <= 0;
        end else if(en) begin
            t12 <= a2;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t13 <= 0;
        end else if(en) begin
            t13 <= b2;
        end
    end
    assign t14 = ($signed(t12) * $signed(t13));
    always @(posedge clock) begin
        if(reset) begin
            t15 <= 0;
        end else if(en) begin
            t15 <= t14;
        end
    end
    assign t16 = ($signed(t15) + $signed(t11));
    always @(posedge clock) begin
        if(reset) begin
            t17 <= 0;
        end else if(en) begin
            t17 <= t16;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t18 <= 0;
        end else if(en) begin
            t18 <= a3;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t19 <= 0;
        end else if(en) begin
            t19 <= b3;
        end
    end
    assign t20 = ($signed(t18) * $signed(t19));
    always @(posedge clock) begin
        if(reset) begin
            t21 <= 0;
        end else if(en) begin
            t21 <= t20;
        end
    end
    assign t22 = ($signed(t21) + $signed(t17));
    always @(posedge clock) begin
        if(reset) begin
            t23 <= 0;
        end else if(en) begin
            t23 <= t22;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t24 <= 0;
        end else if(en) begin
            t24 <= a4;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t25 <= 0;
        end else if(en) begin
            t25 <= b4;
        end
    end
    assign t26 = ($signed(t24) * $signed(t25));
    always @(posedge clock) begin
        if(reset) begin
            t27 <= 0;
        end else if(en) begin
            t27 <= t26;
        end
    end
    assign t28 = ($signed(t27) + $signed(t23));
    always @(posedge clock) begin
        if(reset) begin
            t29 <= 0;
        end else if(en) begin
            t29 <= t28;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t30 <= 0;
        end else if(en) begin
            t30 <= a5;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t31 <= 0;
        end else if(en) begin
            t31 <= b5;
        end
    end
    assign t32 = ($signed(t30) * $signed(t31));
    always @(posedge clock) begin
        if(reset) begin
            t33 <= 0;
        end else if(en) begin
            t33 <= t32;
        end
    end
    assign t34 = ($signed(t33) + $signed(t29));
    always @(posedge clock) begin
        if(reset) begin
            t35 <= 0;
        end else if(en) begin
            t35 <= t34;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t36 <= 0;
        end else if(en) begin
            t36 <= a6;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t37 <= 0;
        end else if(en) begin
            t37 <= b6;
        end
    end
    assign t38 = ($signed(t36) * $signed(t37));
    always @(posedge clock) begin
        if(reset) begin
            t39 <= 0;
        end else if(en) begin
            t39 <= t38;
        end
    end
    assign t40 = ($signed(t39) + $signed(t35));
    always @(posedge clock) begin
        if(reset) begin
            t41 <= 0;
        end else if(en) begin
            t41 <= t40;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t42 <= 0;
        end else if(en) begin
            t42 <= a7;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t43 <= 0;
        end else if(en) begin
            t43 <= b7;
        end
    end
    assign t44 = ($signed(t42) * $signed(t43));
    always @(posedge clock) begin
        if(reset) begin
            t45 <= 0;
        end else if(en) begin
            t45 <= t44;
        end
    end
    assign t46 = ($signed(t45) + $signed(t41));
    always @(posedge clock) begin
        if(reset) begin
            t47 <= 0;
        end else if(en) begin
            t47 <= t46;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t48 <= 0;
        end else if(en) begin
            t48 <= a8;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t49 <= 0;
        end else if(en) begin
            t49 <= b8;
        end
    end
    assign t50 = ($signed(t48) * $signed(t49));
    always @(posedge clock) begin
        if(reset) begin
            t51 <= 0;
        end else if(en) begin
            t51 <= t50;
        end
    end
    assign t52 = ($signed(t51) + $signed(t47));
    always @(posedge clock) begin
        if(reset) begin
            t53 <= 0;
        end else if(en) begin
            t53 <= t52;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t54 <= 0;
        end else if(en) begin
            t54 <= a9;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t55 <= 0;
        end else if(en) begin
            t55 <= b9;
        end
    end
    assign t56 = ($signed(t54) * $signed(t55));
    always @(posedge clock) begin
        if(reset) begin
            t57 <= 0;
        end else if(en) begin
            t57 <= t56;
        end
    end
    assign t58 = ($signed(t57) + $signed(t53));
    always @(posedge clock) begin
        if(reset) begin
            t59 <= 0;
        end else if(en) begin
            t59 <= t58;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t60 <= 0;
        end else if(en) begin
            t60 <= a10;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t61 <= 0;
        end else if(en) begin
            t61 <= b10;
        end
    end
    assign t62 = ($signed(t60) * $signed(t61));
    always @(posedge clock) begin
        if(reset) begin
            t63 <= 0;
        end else if(en) begin
            t63 <= t62;
        end
    end
    assign t64 = ($signed(t63) + $signed(t59));
    always @(posedge clock) begin
        if(reset) begin
            t65 <= 0;
        end else if(en) begin
            t65 <= t64;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t66 <= 0;
        end else if(en) begin
            t66 <= a11;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t67 <= 0;
        end else if(en) begin
            t67 <= b11;
        end
    end
    assign t68 = ($signed(t66) * $signed(t67));
    always @(posedge clock) begin
        if(reset) begin
            t69 <= 0;
        end else if(en) begin
            t69 <= t68;
        end
    end
    assign t70 = ($signed(t69) + $signed(t65));
    always @(posedge clock) begin
        if(reset) begin
            t71 <= 0;
        end else if(en) begin
            t71 <= t70;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t72 <= 0;
        end else if(en) begin
            t72 <= a12;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t73 <= 0;
        end else if(en) begin
            t73 <= b12;
        end
    end
    assign t74 = ($signed(t72) * $signed(t73));
    always @(posedge clock) begin
        if(reset) begin
            t75 <= 0;
        end else if(en) begin
            t75 <= t74;
        end
    end
    assign t76 = ($signed(t75) + $signed(t71));
    always @(posedge clock) begin
        if(reset) begin
            t77 <= 0;
        end else if(en) begin
            t77 <= t76;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t78 <= 0;
        end else if(en) begin
            t78 <= a13;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t79 <= 0;
        end else if(en) begin
            t79 <= b13;
        end
    end
    assign t80 = ($signed(t78) * $signed(t79));
    always @(posedge clock) begin
        if(reset) begin
            t81 <= 0;
        end else if(en) begin
            t81 <= t80;
        end
    end
    assign t82 = ($signed(t81) + $signed(t77));
    always @(posedge clock) begin
        if(reset) begin
            t83 <= 0;
        end else if(en) begin
            t83 <= t82;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t84 <= 0;
        end else if(en) begin
            t84 <= a14;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t85 <= 0;
        end else if(en) begin
            t85 <= b14;
        end
    end
    assign t86 = ($signed(t84) * $signed(t85));
    always @(posedge clock) begin
        if(reset) begin
            t87 <= 0;
        end else if(en) begin
            t87 <= t86;
        end
    end
    assign t88 = ($signed(t87) + $signed(t83));
    always @(posedge clock) begin
        if(reset) begin
            t89 <= 0;
        end else if(en) begin
            t89 <= t88;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t90 <= 0;
        end else if(en) begin
            t90 <= a15;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t91 <= 0;
        end else if(en) begin
            t91 <= b15;
        end
    end
    assign t92 = ($signed(t90) * $signed(t91));
    always @(posedge clock) begin
        if(reset) begin
            t93 <= 0;
        end else if(en) begin
            t93 <= t92;
        end
    end
    assign t94 = ($signed(t93) + $signed(t89));
    always @(posedge clock) begin
        if(reset) begin
            t95 <= 0;
        end else if(en) begin
            t95 <= t94;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t96 <= 0;
        end else if(en) begin
            t96 <= a16;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t97 <= 0;
        end else if(en) begin
            t97 <= b16;
        end
    end
    assign t98 = ($signed(t96) * $signed(t97));
    always @(posedge clock) begin
        if(reset) begin
            t99 <= 0;
        end else if(en) begin
            t99 <= t98;
        end
    end
    assign t100 = ($signed(t99) + $signed(t95));
    always @(posedge clock) begin
        if(reset) begin
            t101 <= 0;
        end else if(en) begin
            t101 <= t100;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t102 <= 0;
        end else if(en) begin
            t102 <= a17;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t103 <= 0;
        end else if(en) begin
            t103 <= b17;
        end
    end
    assign t104 = ($signed(t102) * $signed(t103));
    always @(posedge clock) begin
        if(reset) begin
            t105 <= 0;
        end else if(en) begin
            t105 <= t104;
        end
    end
    assign t106 = ($signed(t105) + $signed(t101));
    always @(posedge clock) begin
        if(reset) begin
            v <= 0;
        end else if(en) begin
            v <= t106;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t108 <= 0;
        end else if(en) begin
            t108 <= c0;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t109 <= 0;
        end else if(en) begin
            t109 <= d0;
        end
    end
    assign t110 = ($signed(t108) * $signed(t109));
    always @(posedge clock) begin
        if(reset) begin
            t111 <= 0;
        end else if(en) begin
            t111 <= t110;
        end
    end
    assign t112 = ($signed(t111) + $signed(n));
    always @(posedge clock) begin
        if(reset) begin
            t113 <= 0;
        end else if(en) begin
            t113 <= t112;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t114 <= 0;
        end else if(en) begin
            t114 <= c1;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t115 <= 0;
        end else if(en) begin
            t115 <= d1;
        end
    end
    assign t116 = ($signed(t114) * $signed(t115));
    always @(posedge clock) begin
        if(reset) begin
            t117 <= 0;
        end else if(en) begin
            t117 <= t116;
        end
    end
    assign t118 = ($signed(t117) + $signed(t113));
    always @(posedge clock) begin
        if(reset) begin
            t119 <= 0;
        end else if(en) begin
            t119 <= t118;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t120 <= 0;
        end else if(en) begin
            t120 <= c2;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t121 <= 0;
        end else if(en) begin
            t121 <= d2;
        end
    end
    assign t122 = ($signed(t120) * $signed(t121));
    always @(posedge clock) begin
        if(reset) begin
            t123 <= 0;
        end else if(en) begin
            t123 <= t122;
        end
    end
    assign t124 = ($signed(t123) + $signed(t119));
    always @(posedge clock) begin
        if(reset) begin
            t125 <= 0;
        end else if(en) begin
            t125 <= t124;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t126 <= 0;
        end else if(en) begin
            t126 <= c3;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t127 <= 0;
        end else if(en) begin
            t127 <= d3;
        end
    end
    assign t128 = ($signed(t126) * $signed(t127));
    always @(posedge clock) begin
        if(reset) begin
            t129 <= 0;
        end else if(en) begin
            t129 <= t128;
        end
    end
    assign t130 = ($signed(t129) + $signed(t125));
    always @(posedge clock) begin
        if(reset) begin
            t131 <= 0;
        end else if(en) begin
            t131 <= t130;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t132 <= 0;
        end else if(en) begin
            t132 <= c4;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t133 <= 0;
        end else if(en) begin
            t133 <= d4;
        end
    end
    assign t134 = ($signed(t132) * $signed(t133));
    always @(posedge clock) begin
        if(reset) begin
            t135 <= 0;
        end else if(en) begin
            t135 <= t134;
        end
    end
    assign t136 = ($signed(t135) + $signed(t131));
    always @(posedge clock) begin
        if(reset) begin
            t137 <= 0;
        end else if(en) begin
            t137 <= t136;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t138 <= 0;
        end else if(en) begin
            t138 <= c5;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t139 <= 0;
        end else if(en) begin
            t139 <= d5;
        end
    end
    assign t140 = ($signed(t138) * $signed(t139));
    always @(posedge clock) begin
        if(reset) begin
            t141 <= 0;
        end else if(en) begin
            t141 <= t140;
        end
    end
    assign t142 = ($signed(t141) + $signed(t137));
    always @(posedge clock) begin
        if(reset) begin
            t143 <= 0;
        end else if(en) begin
            t143 <= t142;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t144 <= 0;
        end else if(en) begin
            t144 <= c6;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t145 <= 0;
        end else if(en) begin
            t145 <= d6;
        end
    end
    assign t146 = ($signed(t144) * $signed(t145));
    always @(posedge clock) begin
        if(reset) begin
            t147 <= 0;
        end else if(en) begin
            t147 <= t146;
        end
    end
    assign t148 = ($signed(t147) + $signed(t143));
    always @(posedge clock) begin
        if(reset) begin
            t149 <= 0;
        end else if(en) begin
            t149 <= t148;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t150 <= 0;
        end else if(en) begin
            t150 <= c7;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t151 <= 0;
        end else if(en) begin
            t151 <= d7;
        end
    end
    assign t152 = ($signed(t150) * $signed(t151));
    always @(posedge clock) begin
        if(reset) begin
            t153 <= 0;
        end else if(en) begin
            t153 <= t152;
        end
    end
    assign t154 = ($signed(t153) + $signed(t149));
    always @(posedge clock) begin
        if(reset) begin
            t155 <= 0;
        end else if(en) begin
            t155 <= t154;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t156 <= 0;
        end else if(en) begin
            t156 <= c8;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t157 <= 0;
        end else if(en) begin
            t157 <= d8;
        end
    end
    assign t158 = ($signed(t156) * $signed(t157));
    always @(posedge clock) begin
        if(reset) begin
            t159 <= 0;
        end else if(en) begin
            t159 <= t158;
        end
    end
    assign t160 = ($signed(t159) + $signed(t155));
    always @(posedge clock) begin
        if(reset) begin
            t161 <= 0;
        end else if(en) begin
            t161 <= t160;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t162 <= 0;
        end else if(en) begin
            t162 <= c9;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t163 <= 0;
        end else if(en) begin
            t163 <= d9;
        end
    end
    assign t164 = ($signed(t162) * $signed(t163));
    always @(posedge clock) begin
        if(reset) begin
            t165 <= 0;
        end else if(en) begin
            t165 <= t164;
        end
    end
    assign t166 = ($signed(t165) + $signed(t161));
    always @(posedge clock) begin
        if(reset) begin
            t167 <= 0;
        end else if(en) begin
            t167 <= t166;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t168 <= 0;
        end else if(en) begin
            t168 <= c10;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t169 <= 0;
        end else if(en) begin
            t169 <= d10;
        end
    end
    assign t170 = ($signed(t168) * $signed(t169));
    always @(posedge clock) begin
        if(reset) begin
            t171 <= 0;
        end else if(en) begin
            t171 <= t170;
        end
    end
    assign t172 = ($signed(t171) + $signed(t167));
    always @(posedge clock) begin
        if(reset) begin
            t173 <= 0;
        end else if(en) begin
            t173 <= t172;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t174 <= 0;
        end else if(en) begin
            t174 <= c11;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t175 <= 0;
        end else if(en) begin
            t175 <= d11;
        end
    end
    assign t176 = ($signed(t174) * $signed(t175));
    always @(posedge clock) begin
        if(reset) begin
            t177 <= 0;
        end else if(en) begin
            t177 <= t176;
        end
    end
    assign t178 = ($signed(t177) + $signed(t173));
    always @(posedge clock) begin
        if(reset) begin
            t179 <= 0;
        end else if(en) begin
            t179 <= t178;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t180 <= 0;
        end else if(en) begin
            t180 <= c12;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t181 <= 0;
        end else if(en) begin
            t181 <= d12;
        end
    end
    assign t182 = ($signed(t180) * $signed(t181));
    always @(posedge clock) begin
        if(reset) begin
            t183 <= 0;
        end else if(en) begin
            t183 <= t182;
        end
    end
    assign t184 = ($signed(t183) + $signed(t179));
    always @(posedge clock) begin
        if(reset) begin
            t185 <= 0;
        end else if(en) begin
            t185 <= t184;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t186 <= 0;
        end else if(en) begin
            t186 <= c13;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t187 <= 0;
        end else if(en) begin
            t187 <= d13;
        end
    end
    assign t188 = ($signed(t186) * $signed(t187));
    always @(posedge clock) begin
        if(reset) begin
            t189 <= 0;
        end else if(en) begin
            t189 <= t188;
        end
    end
    assign t190 = ($signed(t189) + $signed(t185));
    always @(posedge clock) begin
        if(reset) begin
            t191 <= 0;
        end else if(en) begin
            t191 <= t190;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t192 <= 0;
        end else if(en) begin
            t192 <= c14;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t193 <= 0;
        end else if(en) begin
            t193 <= d14;
        end
    end
    assign t194 = ($signed(t192) * $signed(t193));
    always @(posedge clock) begin
        if(reset) begin
            t195 <= 0;
        end else if(en) begin
            t195 <= t194;
        end
    end
    assign t196 = ($signed(t195) + $signed(t191));
    always @(posedge clock) begin
        if(reset) begin
            t197 <= 0;
        end else if(en) begin
            t197 <= t196;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t198 <= 0;
        end else if(en) begin
            t198 <= c15;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t199 <= 0;
        end else if(en) begin
            t199 <= d15;
        end
    end
    assign t200 = ($signed(t198) * $signed(t199));
    always @(posedge clock) begin
        if(reset) begin
            t201 <= 0;
        end else if(en) begin
            t201 <= t200;
        end
    end
    assign t202 = ($signed(t201) + $signed(t197));
    always @(posedge clock) begin
        if(reset) begin
            t203 <= 0;
        end else if(en) begin
            t203 <= t202;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t204 <= 0;
        end else if(en) begin
            t204 <= c16;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t205 <= 0;
        end else if(en) begin
            t205 <= d16;
        end
    end
    assign t206 = ($signed(t204) * $signed(t205));
    always @(posedge clock) begin
        if(reset) begin
            t207 <= 0;
        end else if(en) begin
            t207 <= t206;
        end
    end
    assign t208 = ($signed(t207) + $signed(t203));
    always @(posedge clock) begin
        if(reset) begin
            t209 <= 0;
        end else if(en) begin
            t209 <= t208;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t210 <= 0;
        end else if(en) begin
            t210 <= c17;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t211 <= 0;
        end else if(en) begin
            t211 <= d17;
        end
    end
    assign t212 = ($signed(t210) * $signed(t211));
    always @(posedge clock) begin
        if(reset) begin
            t213 <= 0;
        end else if(en) begin
            t213 <= t212;
        end
    end
    assign t214 = ($signed(t213) + $signed(t209));
    always @(posedge clock) begin
        if(reset) begin
            w <= 0;
        end else if(en) begin
            w <= t214;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t216 <= 0;
        end else if(en) begin
            t216 <= e0;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t217 <= 0;
        end else if(en) begin
            t217 <= f0;
        end
    end
    assign t218 = ($signed(t216) * $signed(t217));
    always @(posedge clock) begin
        if(reset) begin
            t219 <= 0;
        end else if(en) begin
            t219 <= t218;
        end
    end
    assign t220 = ($signed(t219) + $signed(o));
    always @(posedge clock) begin
        if(reset) begin
            t221 <= 0;
        end else if(en) begin
            t221 <= t220;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t222 <= 0;
        end else if(en) begin
            t222 <= e1;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t223 <= 0;
        end else if(en) begin
            t223 <= f1;
        end
    end
    assign t224 = ($signed(t222) * $signed(t223));
    always @(posedge clock) begin
        if(reset) begin
            t225 <= 0;
        end else if(en) begin
            t225 <= t224;
        end
    end
    assign t226 = ($signed(t225) + $signed(t221));
    always @(posedge clock) begin
        if(reset) begin
            t227 <= 0;
        end else if(en) begin
            t227 <= t226;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t228 <= 0;
        end else if(en) begin
            t228 <= e2;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t229 <= 0;
        end else if(en) begin
            t229 <= f2;
        end
    end
    assign t230 = ($signed(t228) * $signed(t229));
    always @(posedge clock) begin
        if(reset) begin
            t231 <= 0;
        end else if(en) begin
            t231 <= t230;
        end
    end
    assign t232 = ($signed(t231) + $signed(t227));
    always @(posedge clock) begin
        if(reset) begin
            t233 <= 0;
        end else if(en) begin
            t233 <= t232;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t234 <= 0;
        end else if(en) begin
            t234 <= e3;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t235 <= 0;
        end else if(en) begin
            t235 <= f3;
        end
    end
    assign t236 = ($signed(t234) * $signed(t235));
    always @(posedge clock) begin
        if(reset) begin
            t237 <= 0;
        end else if(en) begin
            t237 <= t236;
        end
    end
    assign t238 = ($signed(t237) + $signed(t233));
    always @(posedge clock) begin
        if(reset) begin
            t239 <= 0;
        end else if(en) begin
            t239 <= t238;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t240 <= 0;
        end else if(en) begin
            t240 <= e4;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t241 <= 0;
        end else if(en) begin
            t241 <= f4;
        end
    end
    assign t242 = ($signed(t240) * $signed(t241));
    always @(posedge clock) begin
        if(reset) begin
            t243 <= 0;
        end else if(en) begin
            t243 <= t242;
        end
    end
    assign t244 = ($signed(t243) + $signed(t239));
    always @(posedge clock) begin
        if(reset) begin
            t245 <= 0;
        end else if(en) begin
            t245 <= t244;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t246 <= 0;
        end else if(en) begin
            t246 <= e5;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t247 <= 0;
        end else if(en) begin
            t247 <= f5;
        end
    end
    assign t248 = ($signed(t246) * $signed(t247));
    always @(posedge clock) begin
        if(reset) begin
            t249 <= 0;
        end else if(en) begin
            t249 <= t248;
        end
    end
    assign t250 = ($signed(t249) + $signed(t245));
    always @(posedge clock) begin
        if(reset) begin
            t251 <= 0;
        end else if(en) begin
            t251 <= t250;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t252 <= 0;
        end else if(en) begin
            t252 <= e6;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t253 <= 0;
        end else if(en) begin
            t253 <= f6;
        end
    end
    assign t254 = ($signed(t252) * $signed(t253));
    always @(posedge clock) begin
        if(reset) begin
            t255 <= 0;
        end else if(en) begin
            t255 <= t254;
        end
    end
    assign t256 = ($signed(t255) + $signed(t251));
    always @(posedge clock) begin
        if(reset) begin
            t257 <= 0;
        end else if(en) begin
            t257 <= t256;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t258 <= 0;
        end else if(en) begin
            t258 <= e7;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t259 <= 0;
        end else if(en) begin
            t259 <= f7;
        end
    end
    assign t260 = ($signed(t258) * $signed(t259));
    always @(posedge clock) begin
        if(reset) begin
            t261 <= 0;
        end else if(en) begin
            t261 <= t260;
        end
    end
    assign t262 = ($signed(t261) + $signed(t257));
    always @(posedge clock) begin
        if(reset) begin
            t263 <= 0;
        end else if(en) begin
            t263 <= t262;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t264 <= 0;
        end else if(en) begin
            t264 <= e8;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t265 <= 0;
        end else if(en) begin
            t265 <= f8;
        end
    end
    assign t266 = ($signed(t264) * $signed(t265));
    always @(posedge clock) begin
        if(reset) begin
            t267 <= 0;
        end else if(en) begin
            t267 <= t266;
        end
    end
    assign t268 = ($signed(t267) + $signed(t263));
    always @(posedge clock) begin
        if(reset) begin
            t269 <= 0;
        end else if(en) begin
            t269 <= t268;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t270 <= 0;
        end else if(en) begin
            t270 <= e9;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t271 <= 0;
        end else if(en) begin
            t271 <= f9;
        end
    end
    assign t272 = ($signed(t270) * $signed(t271));
    always @(posedge clock) begin
        if(reset) begin
            t273 <= 0;
        end else if(en) begin
            t273 <= t272;
        end
    end
    assign t274 = ($signed(t273) + $signed(t269));
    always @(posedge clock) begin
        if(reset) begin
            t275 <= 0;
        end else if(en) begin
            t275 <= t274;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t276 <= 0;
        end else if(en) begin
            t276 <= e10;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t277 <= 0;
        end else if(en) begin
            t277 <= f10;
        end
    end
    assign t278 = ($signed(t276) * $signed(t277));
    always @(posedge clock) begin
        if(reset) begin
            t279 <= 0;
        end else if(en) begin
            t279 <= t278;
        end
    end
    assign t280 = ($signed(t279) + $signed(t275));
    always @(posedge clock) begin
        if(reset) begin
            t281 <= 0;
        end else if(en) begin
            t281 <= t280;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t282 <= 0;
        end else if(en) begin
            t282 <= e11;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t283 <= 0;
        end else if(en) begin
            t283 <= f11;
        end
    end
    assign t284 = ($signed(t282) * $signed(t283));
    always @(posedge clock) begin
        if(reset) begin
            t285 <= 0;
        end else if(en) begin
            t285 <= t284;
        end
    end
    assign t286 = ($signed(t285) + $signed(t281));
    always @(posedge clock) begin
        if(reset) begin
            t287 <= 0;
        end else if(en) begin
            t287 <= t286;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t288 <= 0;
        end else if(en) begin
            t288 <= e12;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t289 <= 0;
        end else if(en) begin
            t289 <= f12;
        end
    end
    assign t290 = ($signed(t288) * $signed(t289));
    always @(posedge clock) begin
        if(reset) begin
            t291 <= 0;
        end else if(en) begin
            t291 <= t290;
        end
    end
    assign t292 = ($signed(t291) + $signed(t287));
    always @(posedge clock) begin
        if(reset) begin
            t293 <= 0;
        end else if(en) begin
            t293 <= t292;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t294 <= 0;
        end else if(en) begin
            t294 <= e13;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t295 <= 0;
        end else if(en) begin
            t295 <= f13;
        end
    end
    assign t296 = ($signed(t294) * $signed(t295));
    always @(posedge clock) begin
        if(reset) begin
            t297 <= 0;
        end else if(en) begin
            t297 <= t296;
        end
    end
    assign t298 = ($signed(t297) + $signed(t293));
    always @(posedge clock) begin
        if(reset) begin
            t299 <= 0;
        end else if(en) begin
            t299 <= t298;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t300 <= 0;
        end else if(en) begin
            t300 <= e14;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t301 <= 0;
        end else if(en) begin
            t301 <= f14;
        end
    end
    assign t302 = ($signed(t300) * $signed(t301));
    always @(posedge clock) begin
        if(reset) begin
            t303 <= 0;
        end else if(en) begin
            t303 <= t302;
        end
    end
    assign t304 = ($signed(t303) + $signed(t299));
    always @(posedge clock) begin
        if(reset) begin
            t305 <= 0;
        end else if(en) begin
            t305 <= t304;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t306 <= 0;
        end else if(en) begin
            t306 <= e15;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t307 <= 0;
        end else if(en) begin
            t307 <= f15;
        end
    end
    assign t308 = ($signed(t306) * $signed(t307));
    always @(posedge clock) begin
        if(reset) begin
            t309 <= 0;
        end else if(en) begin
            t309 <= t308;
        end
    end
    assign t310 = ($signed(t309) + $signed(t305));
    always @(posedge clock) begin
        if(reset) begin
            t311 <= 0;
        end else if(en) begin
            t311 <= t310;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t312 <= 0;
        end else if(en) begin
            t312 <= e16;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t313 <= 0;
        end else if(en) begin
            t313 <= f16;
        end
    end
    assign t314 = ($signed(t312) * $signed(t313));
    always @(posedge clock) begin
        if(reset) begin
            t315 <= 0;
        end else if(en) begin
            t315 <= t314;
        end
    end
    assign t316 = ($signed(t315) + $signed(t311));
    always @(posedge clock) begin
        if(reset) begin
            t317 <= 0;
        end else if(en) begin
            t317 <= t316;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t318 <= 0;
        end else if(en) begin
            t318 <= e17;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t319 <= 0;
        end else if(en) begin
            t319 <= f17;
        end
    end
    assign t320 = ($signed(t318) * $signed(t319));
    always @(posedge clock) begin
        if(reset) begin
            t321 <= 0;
        end else if(en) begin
            t321 <= t320;
        end
    end
    assign t322 = ($signed(t321) + $signed(t317));
    always @(posedge clock) begin
        if(reset) begin
            x <= 0;
        end else if(en) begin
            x <= t322;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t324 <= 0;
        end else if(en) begin
            t324 <= g0;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t325 <= 0;
        end else if(en) begin
            t325 <= h0;
        end
    end
    assign t326 = ($signed(t324) * $signed(t325));
    always @(posedge clock) begin
        if(reset) begin
            t327 <= 0;
        end else if(en) begin
            t327 <= t326;
        end
    end
    assign t328 = ($signed(t327) + $signed(p));
    always @(posedge clock) begin
        if(reset) begin
            t329 <= 0;
        end else if(en) begin
            t329 <= t328;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t330 <= 0;
        end else if(en) begin
            t330 <= g1;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t331 <= 0;
        end else if(en) begin
            t331 <= h1;
        end
    end
    assign t332 = ($signed(t330) * $signed(t331));
    always @(posedge clock) begin
        if(reset) begin
            t333 <= 0;
        end else if(en) begin
            t333 <= t332;
        end
    end
    assign t334 = ($signed(t333) + $signed(t329));
    always @(posedge clock) begin
        if(reset) begin
            t335 <= 0;
        end else if(en) begin
            t335 <= t334;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t336 <= 0;
        end else if(en) begin
            t336 <= g2;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t337 <= 0;
        end else if(en) begin
            t337 <= h2;
        end
    end
    assign t338 = ($signed(t336) * $signed(t337));
    always @(posedge clock) begin
        if(reset) begin
            t339 <= 0;
        end else if(en) begin
            t339 <= t338;
        end
    end
    assign t340 = ($signed(t339) + $signed(t335));
    always @(posedge clock) begin
        if(reset) begin
            t341 <= 0;
        end else if(en) begin
            t341 <= t340;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t342 <= 0;
        end else if(en) begin
            t342 <= g3;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t343 <= 0;
        end else if(en) begin
            t343 <= h3;
        end
    end
    assign t344 = ($signed(t342) * $signed(t343));
    always @(posedge clock) begin
        if(reset) begin
            t345 <= 0;
        end else if(en) begin
            t345 <= t344;
        end
    end
    assign t346 = ($signed(t345) + $signed(t341));
    always @(posedge clock) begin
        if(reset) begin
            t347 <= 0;
        end else if(en) begin
            t347 <= t346;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t348 <= 0;
        end else if(en) begin
            t348 <= g4;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t349 <= 0;
        end else if(en) begin
            t349 <= h4;
        end
    end
    assign t350 = ($signed(t348) * $signed(t349));
    always @(posedge clock) begin
        if(reset) begin
            t351 <= 0;
        end else if(en) begin
            t351 <= t350;
        end
    end
    assign t352 = ($signed(t351) + $signed(t347));
    always @(posedge clock) begin
        if(reset) begin
            t353 <= 0;
        end else if(en) begin
            t353 <= t352;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t354 <= 0;
        end else if(en) begin
            t354 <= g5;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t355 <= 0;
        end else if(en) begin
            t355 <= h5;
        end
    end
    assign t356 = ($signed(t354) * $signed(t355));
    always @(posedge clock) begin
        if(reset) begin
            t357 <= 0;
        end else if(en) begin
            t357 <= t356;
        end
    end
    assign t358 = ($signed(t357) + $signed(t353));
    always @(posedge clock) begin
        if(reset) begin
            t359 <= 0;
        end else if(en) begin
            t359 <= t358;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t360 <= 0;
        end else if(en) begin
            t360 <= g6;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t361 <= 0;
        end else if(en) begin
            t361 <= h6;
        end
    end
    assign t362 = ($signed(t360) * $signed(t361));
    always @(posedge clock) begin
        if(reset) begin
            t363 <= 0;
        end else if(en) begin
            t363 <= t362;
        end
    end
    assign t364 = ($signed(t363) + $signed(t359));
    always @(posedge clock) begin
        if(reset) begin
            t365 <= 0;
        end else if(en) begin
            t365 <= t364;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t366 <= 0;
        end else if(en) begin
            t366 <= g7;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t367 <= 0;
        end else if(en) begin
            t367 <= h7;
        end
    end
    assign t368 = ($signed(t366) * $signed(t367));
    always @(posedge clock) begin
        if(reset) begin
            t369 <= 0;
        end else if(en) begin
            t369 <= t368;
        end
    end
    assign t370 = ($signed(t369) + $signed(t365));
    always @(posedge clock) begin
        if(reset) begin
            t371 <= 0;
        end else if(en) begin
            t371 <= t370;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t372 <= 0;
        end else if(en) begin
            t372 <= g8;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t373 <= 0;
        end else if(en) begin
            t373 <= h8;
        end
    end
    assign t374 = ($signed(t372) * $signed(t373));
    always @(posedge clock) begin
        if(reset) begin
            t375 <= 0;
        end else if(en) begin
            t375 <= t374;
        end
    end
    assign t376 = ($signed(t375) + $signed(t371));
    always @(posedge clock) begin
        if(reset) begin
            t377 <= 0;
        end else if(en) begin
            t377 <= t376;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t378 <= 0;
        end else if(en) begin
            t378 <= g9;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t379 <= 0;
        end else if(en) begin
            t379 <= h9;
        end
    end
    assign t380 = ($signed(t378) * $signed(t379));
    always @(posedge clock) begin
        if(reset) begin
            t381 <= 0;
        end else if(en) begin
            t381 <= t380;
        end
    end
    assign t382 = ($signed(t381) + $signed(t377));
    always @(posedge clock) begin
        if(reset) begin
            t383 <= 0;
        end else if(en) begin
            t383 <= t382;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t384 <= 0;
        end else if(en) begin
            t384 <= g10;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t385 <= 0;
        end else if(en) begin
            t385 <= h10;
        end
    end
    assign t386 = ($signed(t384) * $signed(t385));
    always @(posedge clock) begin
        if(reset) begin
            t387 <= 0;
        end else if(en) begin
            t387 <= t386;
        end
    end
    assign t388 = ($signed(t387) + $signed(t383));
    always @(posedge clock) begin
        if(reset) begin
            t389 <= 0;
        end else if(en) begin
            t389 <= t388;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t390 <= 0;
        end else if(en) begin
            t390 <= g11;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t391 <= 0;
        end else if(en) begin
            t391 <= h11;
        end
    end
    assign t392 = ($signed(t390) * $signed(t391));
    always @(posedge clock) begin
        if(reset) begin
            t393 <= 0;
        end else if(en) begin
            t393 <= t392;
        end
    end
    assign t394 = ($signed(t393) + $signed(t389));
    always @(posedge clock) begin
        if(reset) begin
            t395 <= 0;
        end else if(en) begin
            t395 <= t394;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t396 <= 0;
        end else if(en) begin
            t396 <= g12;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t397 <= 0;
        end else if(en) begin
            t397 <= h12;
        end
    end
    assign t398 = ($signed(t396) * $signed(t397));
    always @(posedge clock) begin
        if(reset) begin
            t399 <= 0;
        end else if(en) begin
            t399 <= t398;
        end
    end
    assign t400 = ($signed(t399) + $signed(t395));
    always @(posedge clock) begin
        if(reset) begin
            t401 <= 0;
        end else if(en) begin
            t401 <= t400;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t402 <= 0;
        end else if(en) begin
            t402 <= g13;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t403 <= 0;
        end else if(en) begin
            t403 <= h13;
        end
    end
    assign t404 = ($signed(t402) * $signed(t403));
    always @(posedge clock) begin
        if(reset) begin
            t405 <= 0;
        end else if(en) begin
            t405 <= t404;
        end
    end
    assign t406 = ($signed(t405) + $signed(t401));
    always @(posedge clock) begin
        if(reset) begin
            t407 <= 0;
        end else if(en) begin
            t407 <= t406;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t408 <= 0;
        end else if(en) begin
            t408 <= g14;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t409 <= 0;
        end else if(en) begin
            t409 <= h14;
        end
    end
    assign t410 = ($signed(t408) * $signed(t409));
    always @(posedge clock) begin
        if(reset) begin
            t411 <= 0;
        end else if(en) begin
            t411 <= t410;
        end
    end
    assign t412 = ($signed(t411) + $signed(t407));
    always @(posedge clock) begin
        if(reset) begin
            t413 <= 0;
        end else if(en) begin
            t413 <= t412;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t414 <= 0;
        end else if(en) begin
            t414 <= g15;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t415 <= 0;
        end else if(en) begin
            t415 <= h15;
        end
    end
    assign t416 = ($signed(t414) * $signed(t415));
    always @(posedge clock) begin
        if(reset) begin
            t417 <= 0;
        end else if(en) begin
            t417 <= t416;
        end
    end
    assign t418 = ($signed(t417) + $signed(t413));
    always @(posedge clock) begin
        if(reset) begin
            t419 <= 0;
        end else if(en) begin
            t419 <= t418;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t420 <= 0;
        end else if(en) begin
            t420 <= g16;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t421 <= 0;
        end else if(en) begin
            t421 <= h16;
        end
    end
    assign t422 = ($signed(t420) * $signed(t421));
    always @(posedge clock) begin
        if(reset) begin
            t423 <= 0;
        end else if(en) begin
            t423 <= t422;
        end
    end
    assign t424 = ($signed(t423) + $signed(t419));
    always @(posedge clock) begin
        if(reset) begin
            t425 <= 0;
        end else if(en) begin
            t425 <= t424;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t426 <= 0;
        end else if(en) begin
            t426 <= g17;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t427 <= 0;
        end else if(en) begin
            t427 <= h17;
        end
    end
    assign t428 = ($signed(t426) * $signed(t427));
    always @(posedge clock) begin
        if(reset) begin
            t429 <= 0;
        end else if(en) begin
            t429 <= t428;
        end
    end
    assign t430 = ($signed(t429) + $signed(t425));
    always @(posedge clock) begin
        if(reset) begin
            y <= 0;
        end else if(en) begin
            y <= t430;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t432 <= 0;
        end else if(en) begin
            t432 <= i0;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t433 <= 0;
        end else if(en) begin
            t433 <= j0;
        end
    end
    assign t434 = ($signed(t432) * $signed(t433));
    always @(posedge clock) begin
        if(reset) begin
            t435 <= 0;
        end else if(en) begin
            t435 <= t434;
        end
    end
    assign t436 = ($signed(t435) + $signed(q));
    always @(posedge clock) begin
        if(reset) begin
            t437 <= 0;
        end else if(en) begin
            t437 <= t436;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t438 <= 0;
        end else if(en) begin
            t438 <= i1;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t439 <= 0;
        end else if(en) begin
            t439 <= j1;
        end
    end
    assign t440 = ($signed(t438) * $signed(t439));
    always @(posedge clock) begin
        if(reset) begin
            t441 <= 0;
        end else if(en) begin
            t441 <= t440;
        end
    end
    assign t442 = ($signed(t441) + $signed(t437));
    always @(posedge clock) begin
        if(reset) begin
            t443 <= 0;
        end else if(en) begin
            t443 <= t442;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t444 <= 0;
        end else if(en) begin
            t444 <= i2;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t445 <= 0;
        end else if(en) begin
            t445 <= j2;
        end
    end
    assign t446 = ($signed(t444) * $signed(t445));
    always @(posedge clock) begin
        if(reset) begin
            t447 <= 0;
        end else if(en) begin
            t447 <= t446;
        end
    end
    assign t448 = ($signed(t447) + $signed(t443));
    always @(posedge clock) begin
        if(reset) begin
            t449 <= 0;
        end else if(en) begin
            t449 <= t448;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t450 <= 0;
        end else if(en) begin
            t450 <= i3;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t451 <= 0;
        end else if(en) begin
            t451 <= j3;
        end
    end
    assign t452 = ($signed(t450) * $signed(t451));
    always @(posedge clock) begin
        if(reset) begin
            t453 <= 0;
        end else if(en) begin
            t453 <= t452;
        end
    end
    assign t454 = ($signed(t453) + $signed(t449));
    always @(posedge clock) begin
        if(reset) begin
            t455 <= 0;
        end else if(en) begin
            t455 <= t454;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t456 <= 0;
        end else if(en) begin
            t456 <= i4;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t457 <= 0;
        end else if(en) begin
            t457 <= j4;
        end
    end
    assign t458 = ($signed(t456) * $signed(t457));
    always @(posedge clock) begin
        if(reset) begin
            t459 <= 0;
        end else if(en) begin
            t459 <= t458;
        end
    end
    assign t460 = ($signed(t459) + $signed(t455));
    always @(posedge clock) begin
        if(reset) begin
            t461 <= 0;
        end else if(en) begin
            t461 <= t460;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t462 <= 0;
        end else if(en) begin
            t462 <= i5;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t463 <= 0;
        end else if(en) begin
            t463 <= j5;
        end
    end
    assign t464 = ($signed(t462) * $signed(t463));
    always @(posedge clock) begin
        if(reset) begin
            t465 <= 0;
        end else if(en) begin
            t465 <= t464;
        end
    end
    assign t466 = ($signed(t465) + $signed(t461));
    always @(posedge clock) begin
        if(reset) begin
            t467 <= 0;
        end else if(en) begin
            t467 <= t466;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t468 <= 0;
        end else if(en) begin
            t468 <= i6;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t469 <= 0;
        end else if(en) begin
            t469 <= j6;
        end
    end
    assign t470 = ($signed(t468) * $signed(t469));
    always @(posedge clock) begin
        if(reset) begin
            t471 <= 0;
        end else if(en) begin
            t471 <= t470;
        end
    end
    assign t472 = ($signed(t471) + $signed(t467));
    always @(posedge clock) begin
        if(reset) begin
            t473 <= 0;
        end else if(en) begin
            t473 <= t472;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t474 <= 0;
        end else if(en) begin
            t474 <= i7;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t475 <= 0;
        end else if(en) begin
            t475 <= j7;
        end
    end
    assign t476 = ($signed(t474) * $signed(t475));
    always @(posedge clock) begin
        if(reset) begin
            t477 <= 0;
        end else if(en) begin
            t477 <= t476;
        end
    end
    assign t478 = ($signed(t477) + $signed(t473));
    always @(posedge clock) begin
        if(reset) begin
            t479 <= 0;
        end else if(en) begin
            t479 <= t478;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t480 <= 0;
        end else if(en) begin
            t480 <= i8;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t481 <= 0;
        end else if(en) begin
            t481 <= j8;
        end
    end
    assign t482 = ($signed(t480) * $signed(t481));
    always @(posedge clock) begin
        if(reset) begin
            t483 <= 0;
        end else if(en) begin
            t483 <= t482;
        end
    end
    assign t484 = ($signed(t483) + $signed(t479));
    always @(posedge clock) begin
        if(reset) begin
            t485 <= 0;
        end else if(en) begin
            t485 <= t484;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t486 <= 0;
        end else if(en) begin
            t486 <= i9;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t487 <= 0;
        end else if(en) begin
            t487 <= j9;
        end
    end
    assign t488 = ($signed(t486) * $signed(t487));
    always @(posedge clock) begin
        if(reset) begin
            t489 <= 0;
        end else if(en) begin
            t489 <= t488;
        end
    end
    assign t490 = ($signed(t489) + $signed(t485));
    always @(posedge clock) begin
        if(reset) begin
            t491 <= 0;
        end else if(en) begin
            t491 <= t490;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t492 <= 0;
        end else if(en) begin
            t492 <= i10;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t493 <= 0;
        end else if(en) begin
            t493 <= j10;
        end
    end
    assign t494 = ($signed(t492) * $signed(t493));
    always @(posedge clock) begin
        if(reset) begin
            t495 <= 0;
        end else if(en) begin
            t495 <= t494;
        end
    end
    assign t496 = ($signed(t495) + $signed(t491));
    always @(posedge clock) begin
        if(reset) begin
            t497 <= 0;
        end else if(en) begin
            t497 <= t496;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t498 <= 0;
        end else if(en) begin
            t498 <= i11;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t499 <= 0;
        end else if(en) begin
            t499 <= j11;
        end
    end
    assign t500 = ($signed(t498) * $signed(t499));
    always @(posedge clock) begin
        if(reset) begin
            t501 <= 0;
        end else if(en) begin
            t501 <= t500;
        end
    end
    assign t502 = ($signed(t501) + $signed(t497));
    always @(posedge clock) begin
        if(reset) begin
            t503 <= 0;
        end else if(en) begin
            t503 <= t502;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t504 <= 0;
        end else if(en) begin
            t504 <= i12;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t505 <= 0;
        end else if(en) begin
            t505 <= j12;
        end
    end
    assign t506 = ($signed(t504) * $signed(t505));
    always @(posedge clock) begin
        if(reset) begin
            t507 <= 0;
        end else if(en) begin
            t507 <= t506;
        end
    end
    assign t508 = ($signed(t507) + $signed(t503));
    always @(posedge clock) begin
        if(reset) begin
            t509 <= 0;
        end else if(en) begin
            t509 <= t508;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t510 <= 0;
        end else if(en) begin
            t510 <= i13;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t511 <= 0;
        end else if(en) begin
            t511 <= j13;
        end
    end
    assign t512 = ($signed(t510) * $signed(t511));
    always @(posedge clock) begin
        if(reset) begin
            t513 <= 0;
        end else if(en) begin
            t513 <= t512;
        end
    end
    assign t514 = ($signed(t513) + $signed(t509));
    always @(posedge clock) begin
        if(reset) begin
            t515 <= 0;
        end else if(en) begin
            t515 <= t514;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t516 <= 0;
        end else if(en) begin
            t516 <= i14;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t517 <= 0;
        end else if(en) begin
            t517 <= j14;
        end
    end
    assign t518 = ($signed(t516) * $signed(t517));
    always @(posedge clock) begin
        if(reset) begin
            t519 <= 0;
        end else if(en) begin
            t519 <= t518;
        end
    end
    assign t520 = ($signed(t519) + $signed(t515));
    always @(posedge clock) begin
        if(reset) begin
            t521 <= 0;
        end else if(en) begin
            t521 <= t520;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t522 <= 0;
        end else if(en) begin
            t522 <= i15;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t523 <= 0;
        end else if(en) begin
            t523 <= j15;
        end
    end
    assign t524 = ($signed(t522) * $signed(t523));
    always @(posedge clock) begin
        if(reset) begin
            t525 <= 0;
        end else if(en) begin
            t525 <= t524;
        end
    end
    assign t526 = ($signed(t525) + $signed(t521));
    always @(posedge clock) begin
        if(reset) begin
            t527 <= 0;
        end else if(en) begin
            t527 <= t526;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t528 <= 0;
        end else if(en) begin
            t528 <= i16;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t529 <= 0;
        end else if(en) begin
            t529 <= j16;
        end
    end
    assign t530 = ($signed(t528) * $signed(t529));
    always @(posedge clock) begin
        if(reset) begin
            t531 <= 0;
        end else if(en) begin
            t531 <= t530;
        end
    end
    assign t532 = ($signed(t531) + $signed(t527));
    always @(posedge clock) begin
        if(reset) begin
            t533 <= 0;
        end else if(en) begin
            t533 <= t532;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t534 <= 0;
        end else if(en) begin
            t534 <= i17;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t535 <= 0;
        end else if(en) begin
            t535 <= j17;
        end
    end
    assign t536 = ($signed(t534) * $signed(t535));
    always @(posedge clock) begin
        if(reset) begin
            t537 <= 0;
        end else if(en) begin
            t537 <= t536;
        end
    end
    assign t538 = ($signed(t537) + $signed(t533));
    always @(posedge clock) begin
        if(reset) begin
            z <= 0;
        end else if(en) begin
            z <= t538;
        end
    end
endmodule
