module tdot (
    input wire clock,
    input wire reset,
    input wire [7:0] a0,
    input wire [7:0] c0,
    input wire [7:0] e0,
    input wire [7:0] g0,
    input wire [7:0] i0,
    input wire [7:0] a1,
    input wire [7:0] c1,
    input wire [7:0] e1,
    input wire [7:0] g1,
    input wire [7:0] i1,
    input wire [7:0] a2,
    input wire [7:0] c2,
    input wire [7:0] e2,
    input wire [7:0] g2,
    input wire [7:0] i2,
    input wire [7:0] a3,
    input wire [7:0] c3,
    input wire [7:0] e3,
    input wire [7:0] g3,
    input wire [7:0] i3,
    input wire [7:0] a4,
    input wire [7:0] c4,
    input wire [7:0] e4,
    input wire [7:0] g4,
    input wire [7:0] i4,
    input wire [7:0] a5,
    input wire [7:0] c5,
    input wire [7:0] e5,
    input wire [7:0] g5,
    input wire [7:0] i5,
    input wire [7:0] a6,
    input wire [7:0] c6,
    input wire [7:0] e6,
    input wire [7:0] g6,
    input wire [7:0] i6,
    input wire [7:0] a7,
    input wire [7:0] c7,
    input wire [7:0] e7,
    input wire [7:0] g7,
    input wire [7:0] i7,
    input wire [7:0] a8,
    input wire [7:0] c8,
    input wire [7:0] e8,
    input wire [7:0] g8,
    input wire [7:0] i8,
    input wire [7:0] a9,
    input wire [7:0] c9,
    input wire [7:0] e9,
    input wire [7:0] g9,
    input wire [7:0] i9,
    input wire [7:0] a10,
    input wire [7:0] c10,
    input wire [7:0] e10,
    input wire [7:0] g10,
    input wire [7:0] i10,
    input wire [7:0] a11,
    input wire [7:0] c11,
    input wire [7:0] e11,
    input wire [7:0] g11,
    input wire [7:0] i11,
    input wire [7:0] a12,
    input wire [7:0] c12,
    input wire [7:0] e12,
    input wire [7:0] g12,
    input wire [7:0] i12,
    input wire [7:0] a13,
    input wire [7:0] c13,
    input wire [7:0] e13,
    input wire [7:0] g13,
    input wire [7:0] i13,
    input wire [7:0] a14,
    input wire [7:0] c14,
    input wire [7:0] e14,
    input wire [7:0] g14,
    input wire [7:0] i14,
    input wire [7:0] a15,
    input wire [7:0] c15,
    input wire [7:0] e15,
    input wire [7:0] g15,
    input wire [7:0] i15,
    input wire [7:0] a16,
    input wire [7:0] c16,
    input wire [7:0] e16,
    input wire [7:0] g16,
    input wire [7:0] i16,
    input wire [7:0] a17,
    input wire [7:0] c17,
    input wire [7:0] e17,
    input wire [7:0] g17,
    input wire [7:0] i17,
    input wire [7:0] a18,
    input wire [7:0] c18,
    input wire [7:0] e18,
    input wire [7:0] g18,
    input wire [7:0] i18,
    input wire [7:0] a19,
    input wire [7:0] c19,
    input wire [7:0] e19,
    input wire [7:0] g19,
    input wire [7:0] i19,
    input wire [7:0] a20,
    input wire [7:0] c20,
    input wire [7:0] e20,
    input wire [7:0] g20,
    input wire [7:0] i20,
    input wire [7:0] a21,
    input wire [7:0] c21,
    input wire [7:0] e21,
    input wire [7:0] g21,
    input wire [7:0] i21,
    input wire [7:0] a22,
    input wire [7:0] c22,
    input wire [7:0] e22,
    input wire [7:0] g22,
    input wire [7:0] i22,
    input wire [7:0] a23,
    input wire [7:0] c23,
    input wire [7:0] e23,
    input wire [7:0] g23,
    input wire [7:0] i23,
    input wire [7:0] a24,
    input wire [7:0] c24,
    input wire [7:0] e24,
    input wire [7:0] g24,
    input wire [7:0] i24,
    input wire [7:0] a25,
    input wire [7:0] c25,
    input wire [7:0] e25,
    input wire [7:0] g25,
    input wire [7:0] i25,
    input wire [7:0] a26,
    input wire [7:0] c26,
    input wire [7:0] e26,
    input wire [7:0] g26,
    input wire [7:0] i26,
    input wire [7:0] a27,
    input wire [7:0] c27,
    input wire [7:0] e27,
    input wire [7:0] g27,
    input wire [7:0] i27,
    input wire [7:0] a28,
    input wire [7:0] c28,
    input wire [7:0] e28,
    input wire [7:0] g28,
    input wire [7:0] i28,
    input wire [7:0] a29,
    input wire [7:0] c29,
    input wire [7:0] e29,
    input wire [7:0] g29,
    input wire [7:0] i29,
    input wire [7:0] a30,
    input wire [7:0] c30,
    input wire [7:0] e30,
    input wire [7:0] g30,
    input wire [7:0] i30,
    input wire [7:0] a31,
    input wire [7:0] c31,
    input wire [7:0] e31,
    input wire [7:0] g31,
    input wire [7:0] i31,
    input wire [7:0] a32,
    input wire [7:0] c32,
    input wire [7:0] e32,
    input wire [7:0] g32,
    input wire [7:0] i32,
    input wire [7:0] a33,
    input wire [7:0] c33,
    input wire [7:0] e33,
    input wire [7:0] g33,
    input wire [7:0] i33,
    input wire [7:0] a34,
    input wire [7:0] c34,
    input wire [7:0] e34,
    input wire [7:0] g34,
    input wire [7:0] i34,
    input wire [7:0] a35,
    input wire [7:0] c35,
    input wire [7:0] e35,
    input wire [7:0] g35,
    input wire [7:0] i35,
    input wire [7:0] b0,
    input wire [7:0] d0,
    input wire [7:0] f0,
    input wire [7:0] h0,
    input wire [7:0] j0,
    input wire [7:0] b1,
    input wire [7:0] d1,
    input wire [7:0] f1,
    input wire [7:0] h1,
    input wire [7:0] j1,
    input wire [7:0] b2,
    input wire [7:0] d2,
    input wire [7:0] f2,
    input wire [7:0] h2,
    input wire [7:0] j2,
    input wire [7:0] b3,
    input wire [7:0] d3,
    input wire [7:0] f3,
    input wire [7:0] h3,
    input wire [7:0] j3,
    input wire [7:0] b4,
    input wire [7:0] d4,
    input wire [7:0] f4,
    input wire [7:0] h4,
    input wire [7:0] j4,
    input wire [7:0] b5,
    input wire [7:0] d5,
    input wire [7:0] f5,
    input wire [7:0] h5,
    input wire [7:0] j5,
    input wire [7:0] b6,
    input wire [7:0] d6,
    input wire [7:0] f6,
    input wire [7:0] h6,
    input wire [7:0] j6,
    input wire [7:0] b7,
    input wire [7:0] d7,
    input wire [7:0] f7,
    input wire [7:0] h7,
    input wire [7:0] j7,
    input wire [7:0] b8,
    input wire [7:0] d8,
    input wire [7:0] f8,
    input wire [7:0] h8,
    input wire [7:0] j8,
    input wire [7:0] b9,
    input wire [7:0] d9,
    input wire [7:0] f9,
    input wire [7:0] h9,
    input wire [7:0] j9,
    input wire [7:0] b10,
    input wire [7:0] d10,
    input wire [7:0] f10,
    input wire [7:0] h10,
    input wire [7:0] j10,
    input wire [7:0] b11,
    input wire [7:0] d11,
    input wire [7:0] f11,
    input wire [7:0] h11,
    input wire [7:0] j11,
    input wire [7:0] b12,
    input wire [7:0] d12,
    input wire [7:0] f12,
    input wire [7:0] h12,
    input wire [7:0] j12,
    input wire [7:0] b13,
    input wire [7:0] d13,
    input wire [7:0] f13,
    input wire [7:0] h13,
    input wire [7:0] j13,
    input wire [7:0] b14,
    input wire [7:0] d14,
    input wire [7:0] f14,
    input wire [7:0] h14,
    input wire [7:0] j14,
    input wire [7:0] b15,
    input wire [7:0] d15,
    input wire [7:0] f15,
    input wire [7:0] h15,
    input wire [7:0] j15,
    input wire [7:0] b16,
    input wire [7:0] d16,
    input wire [7:0] f16,
    input wire [7:0] h16,
    input wire [7:0] j16,
    input wire [7:0] b17,
    input wire [7:0] d17,
    input wire [7:0] f17,
    input wire [7:0] h17,
    input wire [7:0] j17,
    input wire [7:0] b18,
    input wire [7:0] d18,
    input wire [7:0] f18,
    input wire [7:0] h18,
    input wire [7:0] j18,
    input wire [7:0] b19,
    input wire [7:0] d19,
    input wire [7:0] f19,
    input wire [7:0] h19,
    input wire [7:0] j19,
    input wire [7:0] b20,
    input wire [7:0] d20,
    input wire [7:0] f20,
    input wire [7:0] h20,
    input wire [7:0] j20,
    input wire [7:0] b21,
    input wire [7:0] d21,
    input wire [7:0] f21,
    input wire [7:0] h21,
    input wire [7:0] j21,
    input wire [7:0] b22,
    input wire [7:0] d22,
    input wire [7:0] f22,
    input wire [7:0] h22,
    input wire [7:0] j22,
    input wire [7:0] b23,
    input wire [7:0] d23,
    input wire [7:0] f23,
    input wire [7:0] h23,
    input wire [7:0] j23,
    input wire [7:0] b24,
    input wire [7:0] d24,
    input wire [7:0] f24,
    input wire [7:0] h24,
    input wire [7:0] j24,
    input wire [7:0] b25,
    input wire [7:0] d25,
    input wire [7:0] f25,
    input wire [7:0] h25,
    input wire [7:0] j25,
    input wire [7:0] b26,
    input wire [7:0] d26,
    input wire [7:0] f26,
    input wire [7:0] h26,
    input wire [7:0] j26,
    input wire [7:0] b27,
    input wire [7:0] d27,
    input wire [7:0] f27,
    input wire [7:0] h27,
    input wire [7:0] j27,
    input wire [7:0] b28,
    input wire [7:0] d28,
    input wire [7:0] f28,
    input wire [7:0] h28,
    input wire [7:0] j28,
    input wire [7:0] b29,
    input wire [7:0] d29,
    input wire [7:0] f29,
    input wire [7:0] h29,
    input wire [7:0] j29,
    input wire [7:0] b30,
    input wire [7:0] d30,
    input wire [7:0] f30,
    input wire [7:0] h30,
    input wire [7:0] j30,
    input wire [7:0] b31,
    input wire [7:0] d31,
    input wire [7:0] f31,
    input wire [7:0] h31,
    input wire [7:0] j31,
    input wire [7:0] b32,
    input wire [7:0] d32,
    input wire [7:0] f32,
    input wire [7:0] h32,
    input wire [7:0] j32,
    input wire [7:0] b33,
    input wire [7:0] d33,
    input wire [7:0] f33,
    input wire [7:0] h33,
    input wire [7:0] j33,
    input wire [7:0] b34,
    input wire [7:0] d34,
    input wire [7:0] f34,
    input wire [7:0] h34,
    input wire [7:0] j34,
    input wire [7:0] b35,
    input wire [7:0] d35,
    input wire [7:0] f35,
    input wire [7:0] h35,
    input wire [7:0] j35,
    input wire [7:0] m,
    input wire [7:0] n,
    input wire [7:0] o,
    input wire [7:0] p,
    input wire [7:0] q,
    input wire en,
    output reg [7:0] v,
    output reg [7:0] w,
    output reg [7:0] x,
    output reg [7:0] y,
    output reg [7:0] z
);
    reg [7:0] t0;
    reg [7:0] t1;
    wire [7:0] t2;
    reg [7:0] t3;
    wire [7:0] t4;
    reg [7:0] t5;
    reg [7:0] t6;
    reg [7:0] t7;
    wire [7:0] t8;
    reg [7:0] t9;
    wire [7:0] t10;
    reg [7:0] t11;
    reg [7:0] t12;
    reg [7:0] t13;
    wire [7:0] t14;
    reg [7:0] t15;
    wire [7:0] t16;
    reg [7:0] t17;
    reg [7:0] t18;
    reg [7:0] t19;
    wire [7:0] t20;
    reg [7:0] t21;
    wire [7:0] t22;
    reg [7:0] t23;
    reg [7:0] t24;
    reg [7:0] t25;
    wire [7:0] t26;
    reg [7:0] t27;
    wire [7:0] t28;
    reg [7:0] t29;
    reg [7:0] t30;
    reg [7:0] t31;
    wire [7:0] t32;
    reg [7:0] t33;
    wire [7:0] t34;
    reg [7:0] t35;
    reg [7:0] t36;
    reg [7:0] t37;
    wire [7:0] t38;
    reg [7:0] t39;
    wire [7:0] t40;
    reg [7:0] t41;
    reg [7:0] t42;
    reg [7:0] t43;
    wire [7:0] t44;
    reg [7:0] t45;
    wire [7:0] t46;
    reg [7:0] t47;
    reg [7:0] t48;
    reg [7:0] t49;
    wire [7:0] t50;
    reg [7:0] t51;
    wire [7:0] t52;
    reg [7:0] t53;
    reg [7:0] t54;
    reg [7:0] t55;
    wire [7:0] t56;
    reg [7:0] t57;
    wire [7:0] t58;
    reg [7:0] t59;
    reg [7:0] t60;
    reg [7:0] t61;
    wire [7:0] t62;
    reg [7:0] t63;
    wire [7:0] t64;
    reg [7:0] t65;
    reg [7:0] t66;
    reg [7:0] t67;
    wire [7:0] t68;
    reg [7:0] t69;
    wire [7:0] t70;
    reg [7:0] t71;
    reg [7:0] t72;
    reg [7:0] t73;
    wire [7:0] t74;
    reg [7:0] t75;
    wire [7:0] t76;
    reg [7:0] t77;
    reg [7:0] t78;
    reg [7:0] t79;
    wire [7:0] t80;
    reg [7:0] t81;
    wire [7:0] t82;
    reg [7:0] t83;
    reg [7:0] t84;
    reg [7:0] t85;
    wire [7:0] t86;
    reg [7:0] t87;
    wire [7:0] t88;
    reg [7:0] t89;
    reg [7:0] t90;
    reg [7:0] t91;
    wire [7:0] t92;
    reg [7:0] t93;
    wire [7:0] t94;
    reg [7:0] t95;
    reg [7:0] t96;
    reg [7:0] t97;
    wire [7:0] t98;
    reg [7:0] t99;
    wire [7:0] t100;
    reg [7:0] t101;
    reg [7:0] t102;
    reg [7:0] t103;
    wire [7:0] t104;
    reg [7:0] t105;
    wire [7:0] t106;
    reg [7:0] t107;
    reg [7:0] t108;
    reg [7:0] t109;
    wire [7:0] t110;
    reg [7:0] t111;
    wire [7:0] t112;
    reg [7:0] t113;
    reg [7:0] t114;
    reg [7:0] t115;
    wire [7:0] t116;
    reg [7:0] t117;
    wire [7:0] t118;
    reg [7:0] t119;
    reg [7:0] t120;
    reg [7:0] t121;
    wire [7:0] t122;
    reg [7:0] t123;
    wire [7:0] t124;
    reg [7:0] t125;
    reg [7:0] t126;
    reg [7:0] t127;
    wire [7:0] t128;
    reg [7:0] t129;
    wire [7:0] t130;
    reg [7:0] t131;
    reg [7:0] t132;
    reg [7:0] t133;
    wire [7:0] t134;
    reg [7:0] t135;
    wire [7:0] t136;
    reg [7:0] t137;
    reg [7:0] t138;
    reg [7:0] t139;
    wire [7:0] t140;
    reg [7:0] t141;
    wire [7:0] t142;
    reg [7:0] t143;
    reg [7:0] t144;
    reg [7:0] t145;
    wire [7:0] t146;
    reg [7:0] t147;
    wire [7:0] t148;
    reg [7:0] t149;
    reg [7:0] t150;
    reg [7:0] t151;
    wire [7:0] t152;
    reg [7:0] t153;
    wire [7:0] t154;
    reg [7:0] t155;
    reg [7:0] t156;
    reg [7:0] t157;
    wire [7:0] t158;
    reg [7:0] t159;
    wire [7:0] t160;
    reg [7:0] t161;
    reg [7:0] t162;
    reg [7:0] t163;
    wire [7:0] t164;
    reg [7:0] t165;
    wire [7:0] t166;
    reg [7:0] t167;
    reg [7:0] t168;
    reg [7:0] t169;
    wire [7:0] t170;
    reg [7:0] t171;
    wire [7:0] t172;
    reg [7:0] t173;
    reg [7:0] t174;
    reg [7:0] t175;
    wire [7:0] t176;
    reg [7:0] t177;
    wire [7:0] t178;
    reg [7:0] t179;
    reg [7:0] t180;
    reg [7:0] t181;
    wire [7:0] t182;
    reg [7:0] t183;
    wire [7:0] t184;
    reg [7:0] t185;
    reg [7:0] t186;
    reg [7:0] t187;
    wire [7:0] t188;
    reg [7:0] t189;
    wire [7:0] t190;
    reg [7:0] t191;
    reg [7:0] t192;
    reg [7:0] t193;
    wire [7:0] t194;
    reg [7:0] t195;
    wire [7:0] t196;
    reg [7:0] t197;
    reg [7:0] t198;
    reg [7:0] t199;
    wire [7:0] t200;
    reg [7:0] t201;
    wire [7:0] t202;
    reg [7:0] t203;
    reg [7:0] t204;
    reg [7:0] t205;
    wire [7:0] t206;
    reg [7:0] t207;
    wire [7:0] t208;
    reg [7:0] t209;
    reg [7:0] t210;
    reg [7:0] t211;
    wire [7:0] t212;
    reg [7:0] t213;
    wire [7:0] t214;
    reg [7:0] t216;
    reg [7:0] t217;
    wire [7:0] t218;
    reg [7:0] t219;
    wire [7:0] t220;
    reg [7:0] t221;
    reg [7:0] t222;
    reg [7:0] t223;
    wire [7:0] t224;
    reg [7:0] t225;
    wire [7:0] t226;
    reg [7:0] t227;
    reg [7:0] t228;
    reg [7:0] t229;
    wire [7:0] t230;
    reg [7:0] t231;
    wire [7:0] t232;
    reg [7:0] t233;
    reg [7:0] t234;
    reg [7:0] t235;
    wire [7:0] t236;
    reg [7:0] t237;
    wire [7:0] t238;
    reg [7:0] t239;
    reg [7:0] t240;
    reg [7:0] t241;
    wire [7:0] t242;
    reg [7:0] t243;
    wire [7:0] t244;
    reg [7:0] t245;
    reg [7:0] t246;
    reg [7:0] t247;
    wire [7:0] t248;
    reg [7:0] t249;
    wire [7:0] t250;
    reg [7:0] t251;
    reg [7:0] t252;
    reg [7:0] t253;
    wire [7:0] t254;
    reg [7:0] t255;
    wire [7:0] t256;
    reg [7:0] t257;
    reg [7:0] t258;
    reg [7:0] t259;
    wire [7:0] t260;
    reg [7:0] t261;
    wire [7:0] t262;
    reg [7:0] t263;
    reg [7:0] t264;
    reg [7:0] t265;
    wire [7:0] t266;
    reg [7:0] t267;
    wire [7:0] t268;
    reg [7:0] t269;
    reg [7:0] t270;
    reg [7:0] t271;
    wire [7:0] t272;
    reg [7:0] t273;
    wire [7:0] t274;
    reg [7:0] t275;
    reg [7:0] t276;
    reg [7:0] t277;
    wire [7:0] t278;
    reg [7:0] t279;
    wire [7:0] t280;
    reg [7:0] t281;
    reg [7:0] t282;
    reg [7:0] t283;
    wire [7:0] t284;
    reg [7:0] t285;
    wire [7:0] t286;
    reg [7:0] t287;
    reg [7:0] t288;
    reg [7:0] t289;
    wire [7:0] t290;
    reg [7:0] t291;
    wire [7:0] t292;
    reg [7:0] t293;
    reg [7:0] t294;
    reg [7:0] t295;
    wire [7:0] t296;
    reg [7:0] t297;
    wire [7:0] t298;
    reg [7:0] t299;
    reg [7:0] t300;
    reg [7:0] t301;
    wire [7:0] t302;
    reg [7:0] t303;
    wire [7:0] t304;
    reg [7:0] t305;
    reg [7:0] t306;
    reg [7:0] t307;
    wire [7:0] t308;
    reg [7:0] t309;
    wire [7:0] t310;
    reg [7:0] t311;
    reg [7:0] t312;
    reg [7:0] t313;
    wire [7:0] t314;
    reg [7:0] t315;
    wire [7:0] t316;
    reg [7:0] t317;
    reg [7:0] t318;
    reg [7:0] t319;
    wire [7:0] t320;
    reg [7:0] t321;
    wire [7:0] t322;
    reg [7:0] t323;
    reg [7:0] t324;
    reg [7:0] t325;
    wire [7:0] t326;
    reg [7:0] t327;
    wire [7:0] t328;
    reg [7:0] t329;
    reg [7:0] t330;
    reg [7:0] t331;
    wire [7:0] t332;
    reg [7:0] t333;
    wire [7:0] t334;
    reg [7:0] t335;
    reg [7:0] t336;
    reg [7:0] t337;
    wire [7:0] t338;
    reg [7:0] t339;
    wire [7:0] t340;
    reg [7:0] t341;
    reg [7:0] t342;
    reg [7:0] t343;
    wire [7:0] t344;
    reg [7:0] t345;
    wire [7:0] t346;
    reg [7:0] t347;
    reg [7:0] t348;
    reg [7:0] t349;
    wire [7:0] t350;
    reg [7:0] t351;
    wire [7:0] t352;
    reg [7:0] t353;
    reg [7:0] t354;
    reg [7:0] t355;
    wire [7:0] t356;
    reg [7:0] t357;
    wire [7:0] t358;
    reg [7:0] t359;
    reg [7:0] t360;
    reg [7:0] t361;
    wire [7:0] t362;
    reg [7:0] t363;
    wire [7:0] t364;
    reg [7:0] t365;
    reg [7:0] t366;
    reg [7:0] t367;
    wire [7:0] t368;
    reg [7:0] t369;
    wire [7:0] t370;
    reg [7:0] t371;
    reg [7:0] t372;
    reg [7:0] t373;
    wire [7:0] t374;
    reg [7:0] t375;
    wire [7:0] t376;
    reg [7:0] t377;
    reg [7:0] t378;
    reg [7:0] t379;
    wire [7:0] t380;
    reg [7:0] t381;
    wire [7:0] t382;
    reg [7:0] t383;
    reg [7:0] t384;
    reg [7:0] t385;
    wire [7:0] t386;
    reg [7:0] t387;
    wire [7:0] t388;
    reg [7:0] t389;
    reg [7:0] t390;
    reg [7:0] t391;
    wire [7:0] t392;
    reg [7:0] t393;
    wire [7:0] t394;
    reg [7:0] t395;
    reg [7:0] t396;
    reg [7:0] t397;
    wire [7:0] t398;
    reg [7:0] t399;
    wire [7:0] t400;
    reg [7:0] t401;
    reg [7:0] t402;
    reg [7:0] t403;
    wire [7:0] t404;
    reg [7:0] t405;
    wire [7:0] t406;
    reg [7:0] t407;
    reg [7:0] t408;
    reg [7:0] t409;
    wire [7:0] t410;
    reg [7:0] t411;
    wire [7:0] t412;
    reg [7:0] t413;
    reg [7:0] t414;
    reg [7:0] t415;
    wire [7:0] t416;
    reg [7:0] t417;
    wire [7:0] t418;
    reg [7:0] t419;
    reg [7:0] t420;
    reg [7:0] t421;
    wire [7:0] t422;
    reg [7:0] t423;
    wire [7:0] t424;
    reg [7:0] t425;
    reg [7:0] t426;
    reg [7:0] t427;
    wire [7:0] t428;
    reg [7:0] t429;
    wire [7:0] t430;
    reg [7:0] t432;
    reg [7:0] t433;
    wire [7:0] t434;
    reg [7:0] t435;
    wire [7:0] t436;
    reg [7:0] t437;
    reg [7:0] t438;
    reg [7:0] t439;
    wire [7:0] t440;
    reg [7:0] t441;
    wire [7:0] t442;
    reg [7:0] t443;
    reg [7:0] t444;
    reg [7:0] t445;
    wire [7:0] t446;
    reg [7:0] t447;
    wire [7:0] t448;
    reg [7:0] t449;
    reg [7:0] t450;
    reg [7:0] t451;
    wire [7:0] t452;
    reg [7:0] t453;
    wire [7:0] t454;
    reg [7:0] t455;
    reg [7:0] t456;
    reg [7:0] t457;
    wire [7:0] t458;
    reg [7:0] t459;
    wire [7:0] t460;
    reg [7:0] t461;
    reg [7:0] t462;
    reg [7:0] t463;
    wire [7:0] t464;
    reg [7:0] t465;
    wire [7:0] t466;
    reg [7:0] t467;
    reg [7:0] t468;
    reg [7:0] t469;
    wire [7:0] t470;
    reg [7:0] t471;
    wire [7:0] t472;
    reg [7:0] t473;
    reg [7:0] t474;
    reg [7:0] t475;
    wire [7:0] t476;
    reg [7:0] t477;
    wire [7:0] t478;
    reg [7:0] t479;
    reg [7:0] t480;
    reg [7:0] t481;
    wire [7:0] t482;
    reg [7:0] t483;
    wire [7:0] t484;
    reg [7:0] t485;
    reg [7:0] t486;
    reg [7:0] t487;
    wire [7:0] t488;
    reg [7:0] t489;
    wire [7:0] t490;
    reg [7:0] t491;
    reg [7:0] t492;
    reg [7:0] t493;
    wire [7:0] t494;
    reg [7:0] t495;
    wire [7:0] t496;
    reg [7:0] t497;
    reg [7:0] t498;
    reg [7:0] t499;
    wire [7:0] t500;
    reg [7:0] t501;
    wire [7:0] t502;
    reg [7:0] t503;
    reg [7:0] t504;
    reg [7:0] t505;
    wire [7:0] t506;
    reg [7:0] t507;
    wire [7:0] t508;
    reg [7:0] t509;
    reg [7:0] t510;
    reg [7:0] t511;
    wire [7:0] t512;
    reg [7:0] t513;
    wire [7:0] t514;
    reg [7:0] t515;
    reg [7:0] t516;
    reg [7:0] t517;
    wire [7:0] t518;
    reg [7:0] t519;
    wire [7:0] t520;
    reg [7:0] t521;
    reg [7:0] t522;
    reg [7:0] t523;
    wire [7:0] t524;
    reg [7:0] t525;
    wire [7:0] t526;
    reg [7:0] t527;
    reg [7:0] t528;
    reg [7:0] t529;
    wire [7:0] t530;
    reg [7:0] t531;
    wire [7:0] t532;
    reg [7:0] t533;
    reg [7:0] t534;
    reg [7:0] t535;
    wire [7:0] t536;
    reg [7:0] t537;
    wire [7:0] t538;
    reg [7:0] t539;
    reg [7:0] t540;
    reg [7:0] t541;
    wire [7:0] t542;
    reg [7:0] t543;
    wire [7:0] t544;
    reg [7:0] t545;
    reg [7:0] t546;
    reg [7:0] t547;
    wire [7:0] t548;
    reg [7:0] t549;
    wire [7:0] t550;
    reg [7:0] t551;
    reg [7:0] t552;
    reg [7:0] t553;
    wire [7:0] t554;
    reg [7:0] t555;
    wire [7:0] t556;
    reg [7:0] t557;
    reg [7:0] t558;
    reg [7:0] t559;
    wire [7:0] t560;
    reg [7:0] t561;
    wire [7:0] t562;
    reg [7:0] t563;
    reg [7:0] t564;
    reg [7:0] t565;
    wire [7:0] t566;
    reg [7:0] t567;
    wire [7:0] t568;
    reg [7:0] t569;
    reg [7:0] t570;
    reg [7:0] t571;
    wire [7:0] t572;
    reg [7:0] t573;
    wire [7:0] t574;
    reg [7:0] t575;
    reg [7:0] t576;
    reg [7:0] t577;
    wire [7:0] t578;
    reg [7:0] t579;
    wire [7:0] t580;
    reg [7:0] t581;
    reg [7:0] t582;
    reg [7:0] t583;
    wire [7:0] t584;
    reg [7:0] t585;
    wire [7:0] t586;
    reg [7:0] t587;
    reg [7:0] t588;
    reg [7:0] t589;
    wire [7:0] t590;
    reg [7:0] t591;
    wire [7:0] t592;
    reg [7:0] t593;
    reg [7:0] t594;
    reg [7:0] t595;
    wire [7:0] t596;
    reg [7:0] t597;
    wire [7:0] t598;
    reg [7:0] t599;
    reg [7:0] t600;
    reg [7:0] t601;
    wire [7:0] t602;
    reg [7:0] t603;
    wire [7:0] t604;
    reg [7:0] t605;
    reg [7:0] t606;
    reg [7:0] t607;
    wire [7:0] t608;
    reg [7:0] t609;
    wire [7:0] t610;
    reg [7:0] t611;
    reg [7:0] t612;
    reg [7:0] t613;
    wire [7:0] t614;
    reg [7:0] t615;
    wire [7:0] t616;
    reg [7:0] t617;
    reg [7:0] t618;
    reg [7:0] t619;
    wire [7:0] t620;
    reg [7:0] t621;
    wire [7:0] t622;
    reg [7:0] t623;
    reg [7:0] t624;
    reg [7:0] t625;
    wire [7:0] t626;
    reg [7:0] t627;
    wire [7:0] t628;
    reg [7:0] t629;
    reg [7:0] t630;
    reg [7:0] t631;
    wire [7:0] t632;
    reg [7:0] t633;
    wire [7:0] t634;
    reg [7:0] t635;
    reg [7:0] t636;
    reg [7:0] t637;
    wire [7:0] t638;
    reg [7:0] t639;
    wire [7:0] t640;
    reg [7:0] t641;
    reg [7:0] t642;
    reg [7:0] t643;
    wire [7:0] t644;
    reg [7:0] t645;
    wire [7:0] t646;
    reg [7:0] t648;
    reg [7:0] t649;
    wire [7:0] t650;
    reg [7:0] t651;
    wire [7:0] t652;
    reg [7:0] t653;
    reg [7:0] t654;
    reg [7:0] t655;
    wire [7:0] t656;
    reg [7:0] t657;
    wire [7:0] t658;
    reg [7:0] t659;
    reg [7:0] t660;
    reg [7:0] t661;
    wire [7:0] t662;
    reg [7:0] t663;
    wire [7:0] t664;
    reg [7:0] t665;
    reg [7:0] t666;
    reg [7:0] t667;
    wire [7:0] t668;
    reg [7:0] t669;
    wire [7:0] t670;
    reg [7:0] t671;
    reg [7:0] t672;
    reg [7:0] t673;
    wire [7:0] t674;
    reg [7:0] t675;
    wire [7:0] t676;
    reg [7:0] t677;
    reg [7:0] t678;
    reg [7:0] t679;
    wire [7:0] t680;
    reg [7:0] t681;
    wire [7:0] t682;
    reg [7:0] t683;
    reg [7:0] t684;
    reg [7:0] t685;
    wire [7:0] t686;
    reg [7:0] t687;
    wire [7:0] t688;
    reg [7:0] t689;
    reg [7:0] t690;
    reg [7:0] t691;
    wire [7:0] t692;
    reg [7:0] t693;
    wire [7:0] t694;
    reg [7:0] t695;
    reg [7:0] t696;
    reg [7:0] t697;
    wire [7:0] t698;
    reg [7:0] t699;
    wire [7:0] t700;
    reg [7:0] t701;
    reg [7:0] t702;
    reg [7:0] t703;
    wire [7:0] t704;
    reg [7:0] t705;
    wire [7:0] t706;
    reg [7:0] t707;
    reg [7:0] t708;
    reg [7:0] t709;
    wire [7:0] t710;
    reg [7:0] t711;
    wire [7:0] t712;
    reg [7:0] t713;
    reg [7:0] t714;
    reg [7:0] t715;
    wire [7:0] t716;
    reg [7:0] t717;
    wire [7:0] t718;
    reg [7:0] t719;
    reg [7:0] t720;
    reg [7:0] t721;
    wire [7:0] t722;
    reg [7:0] t723;
    wire [7:0] t724;
    reg [7:0] t725;
    reg [7:0] t726;
    reg [7:0] t727;
    wire [7:0] t728;
    reg [7:0] t729;
    wire [7:0] t730;
    reg [7:0] t731;
    reg [7:0] t732;
    reg [7:0] t733;
    wire [7:0] t734;
    reg [7:0] t735;
    wire [7:0] t736;
    reg [7:0] t737;
    reg [7:0] t738;
    reg [7:0] t739;
    wire [7:0] t740;
    reg [7:0] t741;
    wire [7:0] t742;
    reg [7:0] t743;
    reg [7:0] t744;
    reg [7:0] t745;
    wire [7:0] t746;
    reg [7:0] t747;
    wire [7:0] t748;
    reg [7:0] t749;
    reg [7:0] t750;
    reg [7:0] t751;
    wire [7:0] t752;
    reg [7:0] t753;
    wire [7:0] t754;
    reg [7:0] t755;
    reg [7:0] t756;
    reg [7:0] t757;
    wire [7:0] t758;
    reg [7:0] t759;
    wire [7:0] t760;
    reg [7:0] t761;
    reg [7:0] t762;
    reg [7:0] t763;
    wire [7:0] t764;
    reg [7:0] t765;
    wire [7:0] t766;
    reg [7:0] t767;
    reg [7:0] t768;
    reg [7:0] t769;
    wire [7:0] t770;
    reg [7:0] t771;
    wire [7:0] t772;
    reg [7:0] t773;
    reg [7:0] t774;
    reg [7:0] t775;
    wire [7:0] t776;
    reg [7:0] t777;
    wire [7:0] t778;
    reg [7:0] t779;
    reg [7:0] t780;
    reg [7:0] t781;
    wire [7:0] t782;
    reg [7:0] t783;
    wire [7:0] t784;
    reg [7:0] t785;
    reg [7:0] t786;
    reg [7:0] t787;
    wire [7:0] t788;
    reg [7:0] t789;
    wire [7:0] t790;
    reg [7:0] t791;
    reg [7:0] t792;
    reg [7:0] t793;
    wire [7:0] t794;
    reg [7:0] t795;
    wire [7:0] t796;
    reg [7:0] t797;
    reg [7:0] t798;
    reg [7:0] t799;
    wire [7:0] t800;
    reg [7:0] t801;
    wire [7:0] t802;
    reg [7:0] t803;
    reg [7:0] t804;
    reg [7:0] t805;
    wire [7:0] t806;
    reg [7:0] t807;
    wire [7:0] t808;
    reg [7:0] t809;
    reg [7:0] t810;
    reg [7:0] t811;
    wire [7:0] t812;
    reg [7:0] t813;
    wire [7:0] t814;
    reg [7:0] t815;
    reg [7:0] t816;
    reg [7:0] t817;
    wire [7:0] t818;
    reg [7:0] t819;
    wire [7:0] t820;
    reg [7:0] t821;
    reg [7:0] t822;
    reg [7:0] t823;
    wire [7:0] t824;
    reg [7:0] t825;
    wire [7:0] t826;
    reg [7:0] t827;
    reg [7:0] t828;
    reg [7:0] t829;
    wire [7:0] t830;
    reg [7:0] t831;
    wire [7:0] t832;
    reg [7:0] t833;
    reg [7:0] t834;
    reg [7:0] t835;
    wire [7:0] t836;
    reg [7:0] t837;
    wire [7:0] t838;
    reg [7:0] t839;
    reg [7:0] t840;
    reg [7:0] t841;
    wire [7:0] t842;
    reg [7:0] t843;
    wire [7:0] t844;
    reg [7:0] t845;
    reg [7:0] t846;
    reg [7:0] t847;
    wire [7:0] t848;
    reg [7:0] t849;
    wire [7:0] t850;
    reg [7:0] t851;
    reg [7:0] t852;
    reg [7:0] t853;
    wire [7:0] t854;
    reg [7:0] t855;
    wire [7:0] t856;
    reg [7:0] t857;
    reg [7:0] t858;
    reg [7:0] t859;
    wire [7:0] t860;
    reg [7:0] t861;
    wire [7:0] t862;
    reg [7:0] t864;
    reg [7:0] t865;
    wire [7:0] t866;
    reg [7:0] t867;
    wire [7:0] t868;
    reg [7:0] t869;
    reg [7:0] t870;
    reg [7:0] t871;
    wire [7:0] t872;
    reg [7:0] t873;
    wire [7:0] t874;
    reg [7:0] t875;
    reg [7:0] t876;
    reg [7:0] t877;
    wire [7:0] t878;
    reg [7:0] t879;
    wire [7:0] t880;
    reg [7:0] t881;
    reg [7:0] t882;
    reg [7:0] t883;
    wire [7:0] t884;
    reg [7:0] t885;
    wire [7:0] t886;
    reg [7:0] t887;
    reg [7:0] t888;
    reg [7:0] t889;
    wire [7:0] t890;
    reg [7:0] t891;
    wire [7:0] t892;
    reg [7:0] t893;
    reg [7:0] t894;
    reg [7:0] t895;
    wire [7:0] t896;
    reg [7:0] t897;
    wire [7:0] t898;
    reg [7:0] t899;
    reg [7:0] t900;
    reg [7:0] t901;
    wire [7:0] t902;
    reg [7:0] t903;
    wire [7:0] t904;
    reg [7:0] t905;
    reg [7:0] t906;
    reg [7:0] t907;
    wire [7:0] t908;
    reg [7:0] t909;
    wire [7:0] t910;
    reg [7:0] t911;
    reg [7:0] t912;
    reg [7:0] t913;
    wire [7:0] t914;
    reg [7:0] t915;
    wire [7:0] t916;
    reg [7:0] t917;
    reg [7:0] t918;
    reg [7:0] t919;
    wire [7:0] t920;
    reg [7:0] t921;
    wire [7:0] t922;
    reg [7:0] t923;
    reg [7:0] t924;
    reg [7:0] t925;
    wire [7:0] t926;
    reg [7:0] t927;
    wire [7:0] t928;
    reg [7:0] t929;
    reg [7:0] t930;
    reg [7:0] t931;
    wire [7:0] t932;
    reg [7:0] t933;
    wire [7:0] t934;
    reg [7:0] t935;
    reg [7:0] t936;
    reg [7:0] t937;
    wire [7:0] t938;
    reg [7:0] t939;
    wire [7:0] t940;
    reg [7:0] t941;
    reg [7:0] t942;
    reg [7:0] t943;
    wire [7:0] t944;
    reg [7:0] t945;
    wire [7:0] t946;
    reg [7:0] t947;
    reg [7:0] t948;
    reg [7:0] t949;
    wire [7:0] t950;
    reg [7:0] t951;
    wire [7:0] t952;
    reg [7:0] t953;
    reg [7:0] t954;
    reg [7:0] t955;
    wire [7:0] t956;
    reg [7:0] t957;
    wire [7:0] t958;
    reg [7:0] t959;
    reg [7:0] t960;
    reg [7:0] t961;
    wire [7:0] t962;
    reg [7:0] t963;
    wire [7:0] t964;
    reg [7:0] t965;
    reg [7:0] t966;
    reg [7:0] t967;
    wire [7:0] t968;
    reg [7:0] t969;
    wire [7:0] t970;
    reg [7:0] t971;
    reg [7:0] t972;
    reg [7:0] t973;
    wire [7:0] t974;
    reg [7:0] t975;
    wire [7:0] t976;
    reg [7:0] t977;
    reg [7:0] t978;
    reg [7:0] t979;
    wire [7:0] t980;
    reg [7:0] t981;
    wire [7:0] t982;
    reg [7:0] t983;
    reg [7:0] t984;
    reg [7:0] t985;
    wire [7:0] t986;
    reg [7:0] t987;
    wire [7:0] t988;
    reg [7:0] t989;
    reg [7:0] t990;
    reg [7:0] t991;
    wire [7:0] t992;
    reg [7:0] t993;
    wire [7:0] t994;
    reg [7:0] t995;
    reg [7:0] t996;
    reg [7:0] t997;
    wire [7:0] t998;
    reg [7:0] t999;
    wire [7:0] t1000;
    reg [7:0] t1001;
    reg [7:0] t1002;
    reg [7:0] t1003;
    wire [7:0] t1004;
    reg [7:0] t1005;
    wire [7:0] t1006;
    reg [7:0] t1007;
    reg [7:0] t1008;
    reg [7:0] t1009;
    wire [7:0] t1010;
    reg [7:0] t1011;
    wire [7:0] t1012;
    reg [7:0] t1013;
    reg [7:0] t1014;
    reg [7:0] t1015;
    wire [7:0] t1016;
    reg [7:0] t1017;
    wire [7:0] t1018;
    reg [7:0] t1019;
    reg [7:0] t1020;
    reg [7:0] t1021;
    wire [7:0] t1022;
    reg [7:0] t1023;
    wire [7:0] t1024;
    reg [7:0] t1025;
    reg [7:0] t1026;
    reg [7:0] t1027;
    wire [7:0] t1028;
    reg [7:0] t1029;
    wire [7:0] t1030;
    reg [7:0] t1031;
    reg [7:0] t1032;
    reg [7:0] t1033;
    wire [7:0] t1034;
    reg [7:0] t1035;
    wire [7:0] t1036;
    reg [7:0] t1037;
    reg [7:0] t1038;
    reg [7:0] t1039;
    wire [7:0] t1040;
    reg [7:0] t1041;
    wire [7:0] t1042;
    reg [7:0] t1043;
    reg [7:0] t1044;
    reg [7:0] t1045;
    wire [7:0] t1046;
    reg [7:0] t1047;
    wire [7:0] t1048;
    reg [7:0] t1049;
    reg [7:0] t1050;
    reg [7:0] t1051;
    wire [7:0] t1052;
    reg [7:0] t1053;
    wire [7:0] t1054;
    reg [7:0] t1055;
    reg [7:0] t1056;
    reg [7:0] t1057;
    wire [7:0] t1058;
    reg [7:0] t1059;
    wire [7:0] t1060;
    reg [7:0] t1061;
    reg [7:0] t1062;
    reg [7:0] t1063;
    wire [7:0] t1064;
    reg [7:0] t1065;
    wire [7:0] t1066;
    reg [7:0] t1067;
    reg [7:0] t1068;
    reg [7:0] t1069;
    wire [7:0] t1070;
    reg [7:0] t1071;
    wire [7:0] t1072;
    reg [7:0] t1073;
    reg [7:0] t1074;
    reg [7:0] t1075;
    wire [7:0] t1076;
    reg [7:0] t1077;
    wire [7:0] t1078;
    always @(posedge clock) begin
        if(reset) begin
            t0 <= 0;
        end else if(en) begin
            t0 <= a0;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t1 <= 0;
        end else if(en) begin
            t1 <= b0;
        end
    end
    assign t2 = ($signed(t0) * $signed(t1));
    always @(posedge clock) begin
        if(reset) begin
            t3 <= 0;
        end else if(en) begin
            t3 <= t2;
        end
    end
    assign t4 = ($signed(t3) + $signed(m));
    always @(posedge clock) begin
        if(reset) begin
            t5 <= 0;
        end else if(en) begin
            t5 <= t4;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t6 <= 0;
        end else if(en) begin
            t6 <= a1;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t7 <= 0;
        end else if(en) begin
            t7 <= b1;
        end
    end
    assign t8 = ($signed(t6) * $signed(t7));
    always @(posedge clock) begin
        if(reset) begin
            t9 <= 0;
        end else if(en) begin
            t9 <= t8;
        end
    end
    assign t10 = ($signed(t9) + $signed(t5));
    always @(posedge clock) begin
        if(reset) begin
            t11 <= 0;
        end else if(en) begin
            t11 <= t10;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t12 <= 0;
        end else if(en) begin
            t12 <= a2;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t13 <= 0;
        end else if(en) begin
            t13 <= b2;
        end
    end
    assign t14 = ($signed(t12) * $signed(t13));
    always @(posedge clock) begin
        if(reset) begin
            t15 <= 0;
        end else if(en) begin
            t15 <= t14;
        end
    end
    assign t16 = ($signed(t15) + $signed(t11));
    always @(posedge clock) begin
        if(reset) begin
            t17 <= 0;
        end else if(en) begin
            t17 <= t16;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t18 <= 0;
        end else if(en) begin
            t18 <= a3;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t19 <= 0;
        end else if(en) begin
            t19 <= b3;
        end
    end
    assign t20 = ($signed(t18) * $signed(t19));
    always @(posedge clock) begin
        if(reset) begin
            t21 <= 0;
        end else if(en) begin
            t21 <= t20;
        end
    end
    assign t22 = ($signed(t21) + $signed(t17));
    always @(posedge clock) begin
        if(reset) begin
            t23 <= 0;
        end else if(en) begin
            t23 <= t22;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t24 <= 0;
        end else if(en) begin
            t24 <= a4;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t25 <= 0;
        end else if(en) begin
            t25 <= b4;
        end
    end
    assign t26 = ($signed(t24) * $signed(t25));
    always @(posedge clock) begin
        if(reset) begin
            t27 <= 0;
        end else if(en) begin
            t27 <= t26;
        end
    end
    assign t28 = ($signed(t27) + $signed(t23));
    always @(posedge clock) begin
        if(reset) begin
            t29 <= 0;
        end else if(en) begin
            t29 <= t28;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t30 <= 0;
        end else if(en) begin
            t30 <= a5;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t31 <= 0;
        end else if(en) begin
            t31 <= b5;
        end
    end
    assign t32 = ($signed(t30) * $signed(t31));
    always @(posedge clock) begin
        if(reset) begin
            t33 <= 0;
        end else if(en) begin
            t33 <= t32;
        end
    end
    assign t34 = ($signed(t33) + $signed(t29));
    always @(posedge clock) begin
        if(reset) begin
            t35 <= 0;
        end else if(en) begin
            t35 <= t34;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t36 <= 0;
        end else if(en) begin
            t36 <= a6;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t37 <= 0;
        end else if(en) begin
            t37 <= b6;
        end
    end
    assign t38 = ($signed(t36) * $signed(t37));
    always @(posedge clock) begin
        if(reset) begin
            t39 <= 0;
        end else if(en) begin
            t39 <= t38;
        end
    end
    assign t40 = ($signed(t39) + $signed(t35));
    always @(posedge clock) begin
        if(reset) begin
            t41 <= 0;
        end else if(en) begin
            t41 <= t40;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t42 <= 0;
        end else if(en) begin
            t42 <= a7;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t43 <= 0;
        end else if(en) begin
            t43 <= b7;
        end
    end
    assign t44 = ($signed(t42) * $signed(t43));
    always @(posedge clock) begin
        if(reset) begin
            t45 <= 0;
        end else if(en) begin
            t45 <= t44;
        end
    end
    assign t46 = ($signed(t45) + $signed(t41));
    always @(posedge clock) begin
        if(reset) begin
            t47 <= 0;
        end else if(en) begin
            t47 <= t46;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t48 <= 0;
        end else if(en) begin
            t48 <= a8;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t49 <= 0;
        end else if(en) begin
            t49 <= b8;
        end
    end
    assign t50 = ($signed(t48) * $signed(t49));
    always @(posedge clock) begin
        if(reset) begin
            t51 <= 0;
        end else if(en) begin
            t51 <= t50;
        end
    end
    assign t52 = ($signed(t51) + $signed(t47));
    always @(posedge clock) begin
        if(reset) begin
            t53 <= 0;
        end else if(en) begin
            t53 <= t52;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t54 <= 0;
        end else if(en) begin
            t54 <= a9;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t55 <= 0;
        end else if(en) begin
            t55 <= b9;
        end
    end
    assign t56 = ($signed(t54) * $signed(t55));
    always @(posedge clock) begin
        if(reset) begin
            t57 <= 0;
        end else if(en) begin
            t57 <= t56;
        end
    end
    assign t58 = ($signed(t57) + $signed(t53));
    always @(posedge clock) begin
        if(reset) begin
            t59 <= 0;
        end else if(en) begin
            t59 <= t58;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t60 <= 0;
        end else if(en) begin
            t60 <= a10;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t61 <= 0;
        end else if(en) begin
            t61 <= b10;
        end
    end
    assign t62 = ($signed(t60) * $signed(t61));
    always @(posedge clock) begin
        if(reset) begin
            t63 <= 0;
        end else if(en) begin
            t63 <= t62;
        end
    end
    assign t64 = ($signed(t63) + $signed(t59));
    always @(posedge clock) begin
        if(reset) begin
            t65 <= 0;
        end else if(en) begin
            t65 <= t64;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t66 <= 0;
        end else if(en) begin
            t66 <= a11;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t67 <= 0;
        end else if(en) begin
            t67 <= b11;
        end
    end
    assign t68 = ($signed(t66) * $signed(t67));
    always @(posedge clock) begin
        if(reset) begin
            t69 <= 0;
        end else if(en) begin
            t69 <= t68;
        end
    end
    assign t70 = ($signed(t69) + $signed(t65));
    always @(posedge clock) begin
        if(reset) begin
            t71 <= 0;
        end else if(en) begin
            t71 <= t70;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t72 <= 0;
        end else if(en) begin
            t72 <= a12;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t73 <= 0;
        end else if(en) begin
            t73 <= b12;
        end
    end
    assign t74 = ($signed(t72) * $signed(t73));
    always @(posedge clock) begin
        if(reset) begin
            t75 <= 0;
        end else if(en) begin
            t75 <= t74;
        end
    end
    assign t76 = ($signed(t75) + $signed(t71));
    always @(posedge clock) begin
        if(reset) begin
            t77 <= 0;
        end else if(en) begin
            t77 <= t76;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t78 <= 0;
        end else if(en) begin
            t78 <= a13;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t79 <= 0;
        end else if(en) begin
            t79 <= b13;
        end
    end
    assign t80 = ($signed(t78) * $signed(t79));
    always @(posedge clock) begin
        if(reset) begin
            t81 <= 0;
        end else if(en) begin
            t81 <= t80;
        end
    end
    assign t82 = ($signed(t81) + $signed(t77));
    always @(posedge clock) begin
        if(reset) begin
            t83 <= 0;
        end else if(en) begin
            t83 <= t82;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t84 <= 0;
        end else if(en) begin
            t84 <= a14;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t85 <= 0;
        end else if(en) begin
            t85 <= b14;
        end
    end
    assign t86 = ($signed(t84) * $signed(t85));
    always @(posedge clock) begin
        if(reset) begin
            t87 <= 0;
        end else if(en) begin
            t87 <= t86;
        end
    end
    assign t88 = ($signed(t87) + $signed(t83));
    always @(posedge clock) begin
        if(reset) begin
            t89 <= 0;
        end else if(en) begin
            t89 <= t88;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t90 <= 0;
        end else if(en) begin
            t90 <= a15;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t91 <= 0;
        end else if(en) begin
            t91 <= b15;
        end
    end
    assign t92 = ($signed(t90) * $signed(t91));
    always @(posedge clock) begin
        if(reset) begin
            t93 <= 0;
        end else if(en) begin
            t93 <= t92;
        end
    end
    assign t94 = ($signed(t93) + $signed(t89));
    always @(posedge clock) begin
        if(reset) begin
            t95 <= 0;
        end else if(en) begin
            t95 <= t94;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t96 <= 0;
        end else if(en) begin
            t96 <= a16;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t97 <= 0;
        end else if(en) begin
            t97 <= b16;
        end
    end
    assign t98 = ($signed(t96) * $signed(t97));
    always @(posedge clock) begin
        if(reset) begin
            t99 <= 0;
        end else if(en) begin
            t99 <= t98;
        end
    end
    assign t100 = ($signed(t99) + $signed(t95));
    always @(posedge clock) begin
        if(reset) begin
            t101 <= 0;
        end else if(en) begin
            t101 <= t100;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t102 <= 0;
        end else if(en) begin
            t102 <= a17;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t103 <= 0;
        end else if(en) begin
            t103 <= b17;
        end
    end
    assign t104 = ($signed(t102) * $signed(t103));
    always @(posedge clock) begin
        if(reset) begin
            t105 <= 0;
        end else if(en) begin
            t105 <= t104;
        end
    end
    assign t106 = ($signed(t105) + $signed(t101));
    always @(posedge clock) begin
        if(reset) begin
            t107 <= 0;
        end else if(en) begin
            t107 <= t106;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t108 <= 0;
        end else if(en) begin
            t108 <= a18;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t109 <= 0;
        end else if(en) begin
            t109 <= b18;
        end
    end
    assign t110 = ($signed(t108) * $signed(t109));
    always @(posedge clock) begin
        if(reset) begin
            t111 <= 0;
        end else if(en) begin
            t111 <= t110;
        end
    end
    assign t112 = ($signed(t111) + $signed(t107));
    always @(posedge clock) begin
        if(reset) begin
            t113 <= 0;
        end else if(en) begin
            t113 <= t112;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t114 <= 0;
        end else if(en) begin
            t114 <= a19;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t115 <= 0;
        end else if(en) begin
            t115 <= b19;
        end
    end
    assign t116 = ($signed(t114) * $signed(t115));
    always @(posedge clock) begin
        if(reset) begin
            t117 <= 0;
        end else if(en) begin
            t117 <= t116;
        end
    end
    assign t118 = ($signed(t117) + $signed(t113));
    always @(posedge clock) begin
        if(reset) begin
            t119 <= 0;
        end else if(en) begin
            t119 <= t118;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t120 <= 0;
        end else if(en) begin
            t120 <= a20;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t121 <= 0;
        end else if(en) begin
            t121 <= b20;
        end
    end
    assign t122 = ($signed(t120) * $signed(t121));
    always @(posedge clock) begin
        if(reset) begin
            t123 <= 0;
        end else if(en) begin
            t123 <= t122;
        end
    end
    assign t124 = ($signed(t123) + $signed(t119));
    always @(posedge clock) begin
        if(reset) begin
            t125 <= 0;
        end else if(en) begin
            t125 <= t124;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t126 <= 0;
        end else if(en) begin
            t126 <= a21;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t127 <= 0;
        end else if(en) begin
            t127 <= b21;
        end
    end
    assign t128 = ($signed(t126) * $signed(t127));
    always @(posedge clock) begin
        if(reset) begin
            t129 <= 0;
        end else if(en) begin
            t129 <= t128;
        end
    end
    assign t130 = ($signed(t129) + $signed(t125));
    always @(posedge clock) begin
        if(reset) begin
            t131 <= 0;
        end else if(en) begin
            t131 <= t130;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t132 <= 0;
        end else if(en) begin
            t132 <= a22;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t133 <= 0;
        end else if(en) begin
            t133 <= b22;
        end
    end
    assign t134 = ($signed(t132) * $signed(t133));
    always @(posedge clock) begin
        if(reset) begin
            t135 <= 0;
        end else if(en) begin
            t135 <= t134;
        end
    end
    assign t136 = ($signed(t135) + $signed(t131));
    always @(posedge clock) begin
        if(reset) begin
            t137 <= 0;
        end else if(en) begin
            t137 <= t136;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t138 <= 0;
        end else if(en) begin
            t138 <= a23;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t139 <= 0;
        end else if(en) begin
            t139 <= b23;
        end
    end
    assign t140 = ($signed(t138) * $signed(t139));
    always @(posedge clock) begin
        if(reset) begin
            t141 <= 0;
        end else if(en) begin
            t141 <= t140;
        end
    end
    assign t142 = ($signed(t141) + $signed(t137));
    always @(posedge clock) begin
        if(reset) begin
            t143 <= 0;
        end else if(en) begin
            t143 <= t142;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t144 <= 0;
        end else if(en) begin
            t144 <= a24;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t145 <= 0;
        end else if(en) begin
            t145 <= b24;
        end
    end
    assign t146 = ($signed(t144) * $signed(t145));
    always @(posedge clock) begin
        if(reset) begin
            t147 <= 0;
        end else if(en) begin
            t147 <= t146;
        end
    end
    assign t148 = ($signed(t147) + $signed(t143));
    always @(posedge clock) begin
        if(reset) begin
            t149 <= 0;
        end else if(en) begin
            t149 <= t148;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t150 <= 0;
        end else if(en) begin
            t150 <= a25;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t151 <= 0;
        end else if(en) begin
            t151 <= b25;
        end
    end
    assign t152 = ($signed(t150) * $signed(t151));
    always @(posedge clock) begin
        if(reset) begin
            t153 <= 0;
        end else if(en) begin
            t153 <= t152;
        end
    end
    assign t154 = ($signed(t153) + $signed(t149));
    always @(posedge clock) begin
        if(reset) begin
            t155 <= 0;
        end else if(en) begin
            t155 <= t154;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t156 <= 0;
        end else if(en) begin
            t156 <= a26;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t157 <= 0;
        end else if(en) begin
            t157 <= b26;
        end
    end
    assign t158 = ($signed(t156) * $signed(t157));
    always @(posedge clock) begin
        if(reset) begin
            t159 <= 0;
        end else if(en) begin
            t159 <= t158;
        end
    end
    assign t160 = ($signed(t159) + $signed(t155));
    always @(posedge clock) begin
        if(reset) begin
            t161 <= 0;
        end else if(en) begin
            t161 <= t160;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t162 <= 0;
        end else if(en) begin
            t162 <= a27;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t163 <= 0;
        end else if(en) begin
            t163 <= b27;
        end
    end
    assign t164 = ($signed(t162) * $signed(t163));
    always @(posedge clock) begin
        if(reset) begin
            t165 <= 0;
        end else if(en) begin
            t165 <= t164;
        end
    end
    assign t166 = ($signed(t165) + $signed(t161));
    always @(posedge clock) begin
        if(reset) begin
            t167 <= 0;
        end else if(en) begin
            t167 <= t166;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t168 <= 0;
        end else if(en) begin
            t168 <= a28;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t169 <= 0;
        end else if(en) begin
            t169 <= b28;
        end
    end
    assign t170 = ($signed(t168) * $signed(t169));
    always @(posedge clock) begin
        if(reset) begin
            t171 <= 0;
        end else if(en) begin
            t171 <= t170;
        end
    end
    assign t172 = ($signed(t171) + $signed(t167));
    always @(posedge clock) begin
        if(reset) begin
            t173 <= 0;
        end else if(en) begin
            t173 <= t172;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t174 <= 0;
        end else if(en) begin
            t174 <= a29;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t175 <= 0;
        end else if(en) begin
            t175 <= b29;
        end
    end
    assign t176 = ($signed(t174) * $signed(t175));
    always @(posedge clock) begin
        if(reset) begin
            t177 <= 0;
        end else if(en) begin
            t177 <= t176;
        end
    end
    assign t178 = ($signed(t177) + $signed(t173));
    always @(posedge clock) begin
        if(reset) begin
            t179 <= 0;
        end else if(en) begin
            t179 <= t178;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t180 <= 0;
        end else if(en) begin
            t180 <= a30;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t181 <= 0;
        end else if(en) begin
            t181 <= b30;
        end
    end
    assign t182 = ($signed(t180) * $signed(t181));
    always @(posedge clock) begin
        if(reset) begin
            t183 <= 0;
        end else if(en) begin
            t183 <= t182;
        end
    end
    assign t184 = ($signed(t183) + $signed(t179));
    always @(posedge clock) begin
        if(reset) begin
            t185 <= 0;
        end else if(en) begin
            t185 <= t184;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t186 <= 0;
        end else if(en) begin
            t186 <= a31;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t187 <= 0;
        end else if(en) begin
            t187 <= b31;
        end
    end
    assign t188 = ($signed(t186) * $signed(t187));
    always @(posedge clock) begin
        if(reset) begin
            t189 <= 0;
        end else if(en) begin
            t189 <= t188;
        end
    end
    assign t190 = ($signed(t189) + $signed(t185));
    always @(posedge clock) begin
        if(reset) begin
            t191 <= 0;
        end else if(en) begin
            t191 <= t190;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t192 <= 0;
        end else if(en) begin
            t192 <= a32;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t193 <= 0;
        end else if(en) begin
            t193 <= b32;
        end
    end
    assign t194 = ($signed(t192) * $signed(t193));
    always @(posedge clock) begin
        if(reset) begin
            t195 <= 0;
        end else if(en) begin
            t195 <= t194;
        end
    end
    assign t196 = ($signed(t195) + $signed(t191));
    always @(posedge clock) begin
        if(reset) begin
            t197 <= 0;
        end else if(en) begin
            t197 <= t196;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t198 <= 0;
        end else if(en) begin
            t198 <= a33;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t199 <= 0;
        end else if(en) begin
            t199 <= b33;
        end
    end
    assign t200 = ($signed(t198) * $signed(t199));
    always @(posedge clock) begin
        if(reset) begin
            t201 <= 0;
        end else if(en) begin
            t201 <= t200;
        end
    end
    assign t202 = ($signed(t201) + $signed(t197));
    always @(posedge clock) begin
        if(reset) begin
            t203 <= 0;
        end else if(en) begin
            t203 <= t202;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t204 <= 0;
        end else if(en) begin
            t204 <= a34;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t205 <= 0;
        end else if(en) begin
            t205 <= b34;
        end
    end
    assign t206 = ($signed(t204) * $signed(t205));
    always @(posedge clock) begin
        if(reset) begin
            t207 <= 0;
        end else if(en) begin
            t207 <= t206;
        end
    end
    assign t208 = ($signed(t207) + $signed(t203));
    always @(posedge clock) begin
        if(reset) begin
            t209 <= 0;
        end else if(en) begin
            t209 <= t208;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t210 <= 0;
        end else if(en) begin
            t210 <= a35;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t211 <= 0;
        end else if(en) begin
            t211 <= b35;
        end
    end
    assign t212 = ($signed(t210) * $signed(t211));
    always @(posedge clock) begin
        if(reset) begin
            t213 <= 0;
        end else if(en) begin
            t213 <= t212;
        end
    end
    assign t214 = ($signed(t213) + $signed(t209));
    always @(posedge clock) begin
        if(reset) begin
            v <= 0;
        end else if(en) begin
            v <= t214;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t216 <= 0;
        end else if(en) begin
            t216 <= c0;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t217 <= 0;
        end else if(en) begin
            t217 <= d0;
        end
    end
    assign t218 = ($signed(t216) * $signed(t217));
    always @(posedge clock) begin
        if(reset) begin
            t219 <= 0;
        end else if(en) begin
            t219 <= t218;
        end
    end
    assign t220 = ($signed(t219) + $signed(n));
    always @(posedge clock) begin
        if(reset) begin
            t221 <= 0;
        end else if(en) begin
            t221 <= t220;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t222 <= 0;
        end else if(en) begin
            t222 <= c1;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t223 <= 0;
        end else if(en) begin
            t223 <= d1;
        end
    end
    assign t224 = ($signed(t222) * $signed(t223));
    always @(posedge clock) begin
        if(reset) begin
            t225 <= 0;
        end else if(en) begin
            t225 <= t224;
        end
    end
    assign t226 = ($signed(t225) + $signed(t221));
    always @(posedge clock) begin
        if(reset) begin
            t227 <= 0;
        end else if(en) begin
            t227 <= t226;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t228 <= 0;
        end else if(en) begin
            t228 <= c2;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t229 <= 0;
        end else if(en) begin
            t229 <= d2;
        end
    end
    assign t230 = ($signed(t228) * $signed(t229));
    always @(posedge clock) begin
        if(reset) begin
            t231 <= 0;
        end else if(en) begin
            t231 <= t230;
        end
    end
    assign t232 = ($signed(t231) + $signed(t227));
    always @(posedge clock) begin
        if(reset) begin
            t233 <= 0;
        end else if(en) begin
            t233 <= t232;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t234 <= 0;
        end else if(en) begin
            t234 <= c3;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t235 <= 0;
        end else if(en) begin
            t235 <= d3;
        end
    end
    assign t236 = ($signed(t234) * $signed(t235));
    always @(posedge clock) begin
        if(reset) begin
            t237 <= 0;
        end else if(en) begin
            t237 <= t236;
        end
    end
    assign t238 = ($signed(t237) + $signed(t233));
    always @(posedge clock) begin
        if(reset) begin
            t239 <= 0;
        end else if(en) begin
            t239 <= t238;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t240 <= 0;
        end else if(en) begin
            t240 <= c4;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t241 <= 0;
        end else if(en) begin
            t241 <= d4;
        end
    end
    assign t242 = ($signed(t240) * $signed(t241));
    always @(posedge clock) begin
        if(reset) begin
            t243 <= 0;
        end else if(en) begin
            t243 <= t242;
        end
    end
    assign t244 = ($signed(t243) + $signed(t239));
    always @(posedge clock) begin
        if(reset) begin
            t245 <= 0;
        end else if(en) begin
            t245 <= t244;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t246 <= 0;
        end else if(en) begin
            t246 <= c5;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t247 <= 0;
        end else if(en) begin
            t247 <= d5;
        end
    end
    assign t248 = ($signed(t246) * $signed(t247));
    always @(posedge clock) begin
        if(reset) begin
            t249 <= 0;
        end else if(en) begin
            t249 <= t248;
        end
    end
    assign t250 = ($signed(t249) + $signed(t245));
    always @(posedge clock) begin
        if(reset) begin
            t251 <= 0;
        end else if(en) begin
            t251 <= t250;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t252 <= 0;
        end else if(en) begin
            t252 <= c6;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t253 <= 0;
        end else if(en) begin
            t253 <= d6;
        end
    end
    assign t254 = ($signed(t252) * $signed(t253));
    always @(posedge clock) begin
        if(reset) begin
            t255 <= 0;
        end else if(en) begin
            t255 <= t254;
        end
    end
    assign t256 = ($signed(t255) + $signed(t251));
    always @(posedge clock) begin
        if(reset) begin
            t257 <= 0;
        end else if(en) begin
            t257 <= t256;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t258 <= 0;
        end else if(en) begin
            t258 <= c7;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t259 <= 0;
        end else if(en) begin
            t259 <= d7;
        end
    end
    assign t260 = ($signed(t258) * $signed(t259));
    always @(posedge clock) begin
        if(reset) begin
            t261 <= 0;
        end else if(en) begin
            t261 <= t260;
        end
    end
    assign t262 = ($signed(t261) + $signed(t257));
    always @(posedge clock) begin
        if(reset) begin
            t263 <= 0;
        end else if(en) begin
            t263 <= t262;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t264 <= 0;
        end else if(en) begin
            t264 <= c8;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t265 <= 0;
        end else if(en) begin
            t265 <= d8;
        end
    end
    assign t266 = ($signed(t264) * $signed(t265));
    always @(posedge clock) begin
        if(reset) begin
            t267 <= 0;
        end else if(en) begin
            t267 <= t266;
        end
    end
    assign t268 = ($signed(t267) + $signed(t263));
    always @(posedge clock) begin
        if(reset) begin
            t269 <= 0;
        end else if(en) begin
            t269 <= t268;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t270 <= 0;
        end else if(en) begin
            t270 <= c9;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t271 <= 0;
        end else if(en) begin
            t271 <= d9;
        end
    end
    assign t272 = ($signed(t270) * $signed(t271));
    always @(posedge clock) begin
        if(reset) begin
            t273 <= 0;
        end else if(en) begin
            t273 <= t272;
        end
    end
    assign t274 = ($signed(t273) + $signed(t269));
    always @(posedge clock) begin
        if(reset) begin
            t275 <= 0;
        end else if(en) begin
            t275 <= t274;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t276 <= 0;
        end else if(en) begin
            t276 <= c10;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t277 <= 0;
        end else if(en) begin
            t277 <= d10;
        end
    end
    assign t278 = ($signed(t276) * $signed(t277));
    always @(posedge clock) begin
        if(reset) begin
            t279 <= 0;
        end else if(en) begin
            t279 <= t278;
        end
    end
    assign t280 = ($signed(t279) + $signed(t275));
    always @(posedge clock) begin
        if(reset) begin
            t281 <= 0;
        end else if(en) begin
            t281 <= t280;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t282 <= 0;
        end else if(en) begin
            t282 <= c11;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t283 <= 0;
        end else if(en) begin
            t283 <= d11;
        end
    end
    assign t284 = ($signed(t282) * $signed(t283));
    always @(posedge clock) begin
        if(reset) begin
            t285 <= 0;
        end else if(en) begin
            t285 <= t284;
        end
    end
    assign t286 = ($signed(t285) + $signed(t281));
    always @(posedge clock) begin
        if(reset) begin
            t287 <= 0;
        end else if(en) begin
            t287 <= t286;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t288 <= 0;
        end else if(en) begin
            t288 <= c12;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t289 <= 0;
        end else if(en) begin
            t289 <= d12;
        end
    end
    assign t290 = ($signed(t288) * $signed(t289));
    always @(posedge clock) begin
        if(reset) begin
            t291 <= 0;
        end else if(en) begin
            t291 <= t290;
        end
    end
    assign t292 = ($signed(t291) + $signed(t287));
    always @(posedge clock) begin
        if(reset) begin
            t293 <= 0;
        end else if(en) begin
            t293 <= t292;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t294 <= 0;
        end else if(en) begin
            t294 <= c13;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t295 <= 0;
        end else if(en) begin
            t295 <= d13;
        end
    end
    assign t296 = ($signed(t294) * $signed(t295));
    always @(posedge clock) begin
        if(reset) begin
            t297 <= 0;
        end else if(en) begin
            t297 <= t296;
        end
    end
    assign t298 = ($signed(t297) + $signed(t293));
    always @(posedge clock) begin
        if(reset) begin
            t299 <= 0;
        end else if(en) begin
            t299 <= t298;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t300 <= 0;
        end else if(en) begin
            t300 <= c14;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t301 <= 0;
        end else if(en) begin
            t301 <= d14;
        end
    end
    assign t302 = ($signed(t300) * $signed(t301));
    always @(posedge clock) begin
        if(reset) begin
            t303 <= 0;
        end else if(en) begin
            t303 <= t302;
        end
    end
    assign t304 = ($signed(t303) + $signed(t299));
    always @(posedge clock) begin
        if(reset) begin
            t305 <= 0;
        end else if(en) begin
            t305 <= t304;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t306 <= 0;
        end else if(en) begin
            t306 <= c15;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t307 <= 0;
        end else if(en) begin
            t307 <= d15;
        end
    end
    assign t308 = ($signed(t306) * $signed(t307));
    always @(posedge clock) begin
        if(reset) begin
            t309 <= 0;
        end else if(en) begin
            t309 <= t308;
        end
    end
    assign t310 = ($signed(t309) + $signed(t305));
    always @(posedge clock) begin
        if(reset) begin
            t311 <= 0;
        end else if(en) begin
            t311 <= t310;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t312 <= 0;
        end else if(en) begin
            t312 <= c16;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t313 <= 0;
        end else if(en) begin
            t313 <= d16;
        end
    end
    assign t314 = ($signed(t312) * $signed(t313));
    always @(posedge clock) begin
        if(reset) begin
            t315 <= 0;
        end else if(en) begin
            t315 <= t314;
        end
    end
    assign t316 = ($signed(t315) + $signed(t311));
    always @(posedge clock) begin
        if(reset) begin
            t317 <= 0;
        end else if(en) begin
            t317 <= t316;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t318 <= 0;
        end else if(en) begin
            t318 <= c17;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t319 <= 0;
        end else if(en) begin
            t319 <= d17;
        end
    end
    assign t320 = ($signed(t318) * $signed(t319));
    always @(posedge clock) begin
        if(reset) begin
            t321 <= 0;
        end else if(en) begin
            t321 <= t320;
        end
    end
    assign t322 = ($signed(t321) + $signed(t317));
    always @(posedge clock) begin
        if(reset) begin
            t323 <= 0;
        end else if(en) begin
            t323 <= t322;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t324 <= 0;
        end else if(en) begin
            t324 <= c18;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t325 <= 0;
        end else if(en) begin
            t325 <= d18;
        end
    end
    assign t326 = ($signed(t324) * $signed(t325));
    always @(posedge clock) begin
        if(reset) begin
            t327 <= 0;
        end else if(en) begin
            t327 <= t326;
        end
    end
    assign t328 = ($signed(t327) + $signed(t323));
    always @(posedge clock) begin
        if(reset) begin
            t329 <= 0;
        end else if(en) begin
            t329 <= t328;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t330 <= 0;
        end else if(en) begin
            t330 <= c19;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t331 <= 0;
        end else if(en) begin
            t331 <= d19;
        end
    end
    assign t332 = ($signed(t330) * $signed(t331));
    always @(posedge clock) begin
        if(reset) begin
            t333 <= 0;
        end else if(en) begin
            t333 <= t332;
        end
    end
    assign t334 = ($signed(t333) + $signed(t329));
    always @(posedge clock) begin
        if(reset) begin
            t335 <= 0;
        end else if(en) begin
            t335 <= t334;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t336 <= 0;
        end else if(en) begin
            t336 <= c20;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t337 <= 0;
        end else if(en) begin
            t337 <= d20;
        end
    end
    assign t338 = ($signed(t336) * $signed(t337));
    always @(posedge clock) begin
        if(reset) begin
            t339 <= 0;
        end else if(en) begin
            t339 <= t338;
        end
    end
    assign t340 = ($signed(t339) + $signed(t335));
    always @(posedge clock) begin
        if(reset) begin
            t341 <= 0;
        end else if(en) begin
            t341 <= t340;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t342 <= 0;
        end else if(en) begin
            t342 <= c21;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t343 <= 0;
        end else if(en) begin
            t343 <= d21;
        end
    end
    assign t344 = ($signed(t342) * $signed(t343));
    always @(posedge clock) begin
        if(reset) begin
            t345 <= 0;
        end else if(en) begin
            t345 <= t344;
        end
    end
    assign t346 = ($signed(t345) + $signed(t341));
    always @(posedge clock) begin
        if(reset) begin
            t347 <= 0;
        end else if(en) begin
            t347 <= t346;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t348 <= 0;
        end else if(en) begin
            t348 <= c22;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t349 <= 0;
        end else if(en) begin
            t349 <= d22;
        end
    end
    assign t350 = ($signed(t348) * $signed(t349));
    always @(posedge clock) begin
        if(reset) begin
            t351 <= 0;
        end else if(en) begin
            t351 <= t350;
        end
    end
    assign t352 = ($signed(t351) + $signed(t347));
    always @(posedge clock) begin
        if(reset) begin
            t353 <= 0;
        end else if(en) begin
            t353 <= t352;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t354 <= 0;
        end else if(en) begin
            t354 <= c23;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t355 <= 0;
        end else if(en) begin
            t355 <= d23;
        end
    end
    assign t356 = ($signed(t354) * $signed(t355));
    always @(posedge clock) begin
        if(reset) begin
            t357 <= 0;
        end else if(en) begin
            t357 <= t356;
        end
    end
    assign t358 = ($signed(t357) + $signed(t353));
    always @(posedge clock) begin
        if(reset) begin
            t359 <= 0;
        end else if(en) begin
            t359 <= t358;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t360 <= 0;
        end else if(en) begin
            t360 <= c24;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t361 <= 0;
        end else if(en) begin
            t361 <= d24;
        end
    end
    assign t362 = ($signed(t360) * $signed(t361));
    always @(posedge clock) begin
        if(reset) begin
            t363 <= 0;
        end else if(en) begin
            t363 <= t362;
        end
    end
    assign t364 = ($signed(t363) + $signed(t359));
    always @(posedge clock) begin
        if(reset) begin
            t365 <= 0;
        end else if(en) begin
            t365 <= t364;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t366 <= 0;
        end else if(en) begin
            t366 <= c25;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t367 <= 0;
        end else if(en) begin
            t367 <= d25;
        end
    end
    assign t368 = ($signed(t366) * $signed(t367));
    always @(posedge clock) begin
        if(reset) begin
            t369 <= 0;
        end else if(en) begin
            t369 <= t368;
        end
    end
    assign t370 = ($signed(t369) + $signed(t365));
    always @(posedge clock) begin
        if(reset) begin
            t371 <= 0;
        end else if(en) begin
            t371 <= t370;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t372 <= 0;
        end else if(en) begin
            t372 <= c26;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t373 <= 0;
        end else if(en) begin
            t373 <= d26;
        end
    end
    assign t374 = ($signed(t372) * $signed(t373));
    always @(posedge clock) begin
        if(reset) begin
            t375 <= 0;
        end else if(en) begin
            t375 <= t374;
        end
    end
    assign t376 = ($signed(t375) + $signed(t371));
    always @(posedge clock) begin
        if(reset) begin
            t377 <= 0;
        end else if(en) begin
            t377 <= t376;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t378 <= 0;
        end else if(en) begin
            t378 <= c27;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t379 <= 0;
        end else if(en) begin
            t379 <= d27;
        end
    end
    assign t380 = ($signed(t378) * $signed(t379));
    always @(posedge clock) begin
        if(reset) begin
            t381 <= 0;
        end else if(en) begin
            t381 <= t380;
        end
    end
    assign t382 = ($signed(t381) + $signed(t377));
    always @(posedge clock) begin
        if(reset) begin
            t383 <= 0;
        end else if(en) begin
            t383 <= t382;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t384 <= 0;
        end else if(en) begin
            t384 <= c28;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t385 <= 0;
        end else if(en) begin
            t385 <= d28;
        end
    end
    assign t386 = ($signed(t384) * $signed(t385));
    always @(posedge clock) begin
        if(reset) begin
            t387 <= 0;
        end else if(en) begin
            t387 <= t386;
        end
    end
    assign t388 = ($signed(t387) + $signed(t383));
    always @(posedge clock) begin
        if(reset) begin
            t389 <= 0;
        end else if(en) begin
            t389 <= t388;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t390 <= 0;
        end else if(en) begin
            t390 <= c29;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t391 <= 0;
        end else if(en) begin
            t391 <= d29;
        end
    end
    assign t392 = ($signed(t390) * $signed(t391));
    always @(posedge clock) begin
        if(reset) begin
            t393 <= 0;
        end else if(en) begin
            t393 <= t392;
        end
    end
    assign t394 = ($signed(t393) + $signed(t389));
    always @(posedge clock) begin
        if(reset) begin
            t395 <= 0;
        end else if(en) begin
            t395 <= t394;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t396 <= 0;
        end else if(en) begin
            t396 <= c30;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t397 <= 0;
        end else if(en) begin
            t397 <= d30;
        end
    end
    assign t398 = ($signed(t396) * $signed(t397));
    always @(posedge clock) begin
        if(reset) begin
            t399 <= 0;
        end else if(en) begin
            t399 <= t398;
        end
    end
    assign t400 = ($signed(t399) + $signed(t395));
    always @(posedge clock) begin
        if(reset) begin
            t401 <= 0;
        end else if(en) begin
            t401 <= t400;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t402 <= 0;
        end else if(en) begin
            t402 <= c31;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t403 <= 0;
        end else if(en) begin
            t403 <= d31;
        end
    end
    assign t404 = ($signed(t402) * $signed(t403));
    always @(posedge clock) begin
        if(reset) begin
            t405 <= 0;
        end else if(en) begin
            t405 <= t404;
        end
    end
    assign t406 = ($signed(t405) + $signed(t401));
    always @(posedge clock) begin
        if(reset) begin
            t407 <= 0;
        end else if(en) begin
            t407 <= t406;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t408 <= 0;
        end else if(en) begin
            t408 <= c32;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t409 <= 0;
        end else if(en) begin
            t409 <= d32;
        end
    end
    assign t410 = ($signed(t408) * $signed(t409));
    always @(posedge clock) begin
        if(reset) begin
            t411 <= 0;
        end else if(en) begin
            t411 <= t410;
        end
    end
    assign t412 = ($signed(t411) + $signed(t407));
    always @(posedge clock) begin
        if(reset) begin
            t413 <= 0;
        end else if(en) begin
            t413 <= t412;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t414 <= 0;
        end else if(en) begin
            t414 <= c33;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t415 <= 0;
        end else if(en) begin
            t415 <= d33;
        end
    end
    assign t416 = ($signed(t414) * $signed(t415));
    always @(posedge clock) begin
        if(reset) begin
            t417 <= 0;
        end else if(en) begin
            t417 <= t416;
        end
    end
    assign t418 = ($signed(t417) + $signed(t413));
    always @(posedge clock) begin
        if(reset) begin
            t419 <= 0;
        end else if(en) begin
            t419 <= t418;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t420 <= 0;
        end else if(en) begin
            t420 <= c34;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t421 <= 0;
        end else if(en) begin
            t421 <= d34;
        end
    end
    assign t422 = ($signed(t420) * $signed(t421));
    always @(posedge clock) begin
        if(reset) begin
            t423 <= 0;
        end else if(en) begin
            t423 <= t422;
        end
    end
    assign t424 = ($signed(t423) + $signed(t419));
    always @(posedge clock) begin
        if(reset) begin
            t425 <= 0;
        end else if(en) begin
            t425 <= t424;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t426 <= 0;
        end else if(en) begin
            t426 <= c35;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t427 <= 0;
        end else if(en) begin
            t427 <= d35;
        end
    end
    assign t428 = ($signed(t426) * $signed(t427));
    always @(posedge clock) begin
        if(reset) begin
            t429 <= 0;
        end else if(en) begin
            t429 <= t428;
        end
    end
    assign t430 = ($signed(t429) + $signed(t425));
    always @(posedge clock) begin
        if(reset) begin
            w <= 0;
        end else if(en) begin
            w <= t430;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t432 <= 0;
        end else if(en) begin
            t432 <= e0;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t433 <= 0;
        end else if(en) begin
            t433 <= f0;
        end
    end
    assign t434 = ($signed(t432) * $signed(t433));
    always @(posedge clock) begin
        if(reset) begin
            t435 <= 0;
        end else if(en) begin
            t435 <= t434;
        end
    end
    assign t436 = ($signed(t435) + $signed(o));
    always @(posedge clock) begin
        if(reset) begin
            t437 <= 0;
        end else if(en) begin
            t437 <= t436;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t438 <= 0;
        end else if(en) begin
            t438 <= e1;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t439 <= 0;
        end else if(en) begin
            t439 <= f1;
        end
    end
    assign t440 = ($signed(t438) * $signed(t439));
    always @(posedge clock) begin
        if(reset) begin
            t441 <= 0;
        end else if(en) begin
            t441 <= t440;
        end
    end
    assign t442 = ($signed(t441) + $signed(t437));
    always @(posedge clock) begin
        if(reset) begin
            t443 <= 0;
        end else if(en) begin
            t443 <= t442;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t444 <= 0;
        end else if(en) begin
            t444 <= e2;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t445 <= 0;
        end else if(en) begin
            t445 <= f2;
        end
    end
    assign t446 = ($signed(t444) * $signed(t445));
    always @(posedge clock) begin
        if(reset) begin
            t447 <= 0;
        end else if(en) begin
            t447 <= t446;
        end
    end
    assign t448 = ($signed(t447) + $signed(t443));
    always @(posedge clock) begin
        if(reset) begin
            t449 <= 0;
        end else if(en) begin
            t449 <= t448;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t450 <= 0;
        end else if(en) begin
            t450 <= e3;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t451 <= 0;
        end else if(en) begin
            t451 <= f3;
        end
    end
    assign t452 = ($signed(t450) * $signed(t451));
    always @(posedge clock) begin
        if(reset) begin
            t453 <= 0;
        end else if(en) begin
            t453 <= t452;
        end
    end
    assign t454 = ($signed(t453) + $signed(t449));
    always @(posedge clock) begin
        if(reset) begin
            t455 <= 0;
        end else if(en) begin
            t455 <= t454;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t456 <= 0;
        end else if(en) begin
            t456 <= e4;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t457 <= 0;
        end else if(en) begin
            t457 <= f4;
        end
    end
    assign t458 = ($signed(t456) * $signed(t457));
    always @(posedge clock) begin
        if(reset) begin
            t459 <= 0;
        end else if(en) begin
            t459 <= t458;
        end
    end
    assign t460 = ($signed(t459) + $signed(t455));
    always @(posedge clock) begin
        if(reset) begin
            t461 <= 0;
        end else if(en) begin
            t461 <= t460;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t462 <= 0;
        end else if(en) begin
            t462 <= e5;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t463 <= 0;
        end else if(en) begin
            t463 <= f5;
        end
    end
    assign t464 = ($signed(t462) * $signed(t463));
    always @(posedge clock) begin
        if(reset) begin
            t465 <= 0;
        end else if(en) begin
            t465 <= t464;
        end
    end
    assign t466 = ($signed(t465) + $signed(t461));
    always @(posedge clock) begin
        if(reset) begin
            t467 <= 0;
        end else if(en) begin
            t467 <= t466;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t468 <= 0;
        end else if(en) begin
            t468 <= e6;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t469 <= 0;
        end else if(en) begin
            t469 <= f6;
        end
    end
    assign t470 = ($signed(t468) * $signed(t469));
    always @(posedge clock) begin
        if(reset) begin
            t471 <= 0;
        end else if(en) begin
            t471 <= t470;
        end
    end
    assign t472 = ($signed(t471) + $signed(t467));
    always @(posedge clock) begin
        if(reset) begin
            t473 <= 0;
        end else if(en) begin
            t473 <= t472;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t474 <= 0;
        end else if(en) begin
            t474 <= e7;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t475 <= 0;
        end else if(en) begin
            t475 <= f7;
        end
    end
    assign t476 = ($signed(t474) * $signed(t475));
    always @(posedge clock) begin
        if(reset) begin
            t477 <= 0;
        end else if(en) begin
            t477 <= t476;
        end
    end
    assign t478 = ($signed(t477) + $signed(t473));
    always @(posedge clock) begin
        if(reset) begin
            t479 <= 0;
        end else if(en) begin
            t479 <= t478;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t480 <= 0;
        end else if(en) begin
            t480 <= e8;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t481 <= 0;
        end else if(en) begin
            t481 <= f8;
        end
    end
    assign t482 = ($signed(t480) * $signed(t481));
    always @(posedge clock) begin
        if(reset) begin
            t483 <= 0;
        end else if(en) begin
            t483 <= t482;
        end
    end
    assign t484 = ($signed(t483) + $signed(t479));
    always @(posedge clock) begin
        if(reset) begin
            t485 <= 0;
        end else if(en) begin
            t485 <= t484;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t486 <= 0;
        end else if(en) begin
            t486 <= e9;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t487 <= 0;
        end else if(en) begin
            t487 <= f9;
        end
    end
    assign t488 = ($signed(t486) * $signed(t487));
    always @(posedge clock) begin
        if(reset) begin
            t489 <= 0;
        end else if(en) begin
            t489 <= t488;
        end
    end
    assign t490 = ($signed(t489) + $signed(t485));
    always @(posedge clock) begin
        if(reset) begin
            t491 <= 0;
        end else if(en) begin
            t491 <= t490;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t492 <= 0;
        end else if(en) begin
            t492 <= e10;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t493 <= 0;
        end else if(en) begin
            t493 <= f10;
        end
    end
    assign t494 = ($signed(t492) * $signed(t493));
    always @(posedge clock) begin
        if(reset) begin
            t495 <= 0;
        end else if(en) begin
            t495 <= t494;
        end
    end
    assign t496 = ($signed(t495) + $signed(t491));
    always @(posedge clock) begin
        if(reset) begin
            t497 <= 0;
        end else if(en) begin
            t497 <= t496;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t498 <= 0;
        end else if(en) begin
            t498 <= e11;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t499 <= 0;
        end else if(en) begin
            t499 <= f11;
        end
    end
    assign t500 = ($signed(t498) * $signed(t499));
    always @(posedge clock) begin
        if(reset) begin
            t501 <= 0;
        end else if(en) begin
            t501 <= t500;
        end
    end
    assign t502 = ($signed(t501) + $signed(t497));
    always @(posedge clock) begin
        if(reset) begin
            t503 <= 0;
        end else if(en) begin
            t503 <= t502;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t504 <= 0;
        end else if(en) begin
            t504 <= e12;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t505 <= 0;
        end else if(en) begin
            t505 <= f12;
        end
    end
    assign t506 = ($signed(t504) * $signed(t505));
    always @(posedge clock) begin
        if(reset) begin
            t507 <= 0;
        end else if(en) begin
            t507 <= t506;
        end
    end
    assign t508 = ($signed(t507) + $signed(t503));
    always @(posedge clock) begin
        if(reset) begin
            t509 <= 0;
        end else if(en) begin
            t509 <= t508;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t510 <= 0;
        end else if(en) begin
            t510 <= e13;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t511 <= 0;
        end else if(en) begin
            t511 <= f13;
        end
    end
    assign t512 = ($signed(t510) * $signed(t511));
    always @(posedge clock) begin
        if(reset) begin
            t513 <= 0;
        end else if(en) begin
            t513 <= t512;
        end
    end
    assign t514 = ($signed(t513) + $signed(t509));
    always @(posedge clock) begin
        if(reset) begin
            t515 <= 0;
        end else if(en) begin
            t515 <= t514;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t516 <= 0;
        end else if(en) begin
            t516 <= e14;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t517 <= 0;
        end else if(en) begin
            t517 <= f14;
        end
    end
    assign t518 = ($signed(t516) * $signed(t517));
    always @(posedge clock) begin
        if(reset) begin
            t519 <= 0;
        end else if(en) begin
            t519 <= t518;
        end
    end
    assign t520 = ($signed(t519) + $signed(t515));
    always @(posedge clock) begin
        if(reset) begin
            t521 <= 0;
        end else if(en) begin
            t521 <= t520;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t522 <= 0;
        end else if(en) begin
            t522 <= e15;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t523 <= 0;
        end else if(en) begin
            t523 <= f15;
        end
    end
    assign t524 = ($signed(t522) * $signed(t523));
    always @(posedge clock) begin
        if(reset) begin
            t525 <= 0;
        end else if(en) begin
            t525 <= t524;
        end
    end
    assign t526 = ($signed(t525) + $signed(t521));
    always @(posedge clock) begin
        if(reset) begin
            t527 <= 0;
        end else if(en) begin
            t527 <= t526;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t528 <= 0;
        end else if(en) begin
            t528 <= e16;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t529 <= 0;
        end else if(en) begin
            t529 <= f16;
        end
    end
    assign t530 = ($signed(t528) * $signed(t529));
    always @(posedge clock) begin
        if(reset) begin
            t531 <= 0;
        end else if(en) begin
            t531 <= t530;
        end
    end
    assign t532 = ($signed(t531) + $signed(t527));
    always @(posedge clock) begin
        if(reset) begin
            t533 <= 0;
        end else if(en) begin
            t533 <= t532;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t534 <= 0;
        end else if(en) begin
            t534 <= e17;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t535 <= 0;
        end else if(en) begin
            t535 <= f17;
        end
    end
    assign t536 = ($signed(t534) * $signed(t535));
    always @(posedge clock) begin
        if(reset) begin
            t537 <= 0;
        end else if(en) begin
            t537 <= t536;
        end
    end
    assign t538 = ($signed(t537) + $signed(t533));
    always @(posedge clock) begin
        if(reset) begin
            t539 <= 0;
        end else if(en) begin
            t539 <= t538;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t540 <= 0;
        end else if(en) begin
            t540 <= e18;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t541 <= 0;
        end else if(en) begin
            t541 <= f18;
        end
    end
    assign t542 = ($signed(t540) * $signed(t541));
    always @(posedge clock) begin
        if(reset) begin
            t543 <= 0;
        end else if(en) begin
            t543 <= t542;
        end
    end
    assign t544 = ($signed(t543) + $signed(t539));
    always @(posedge clock) begin
        if(reset) begin
            t545 <= 0;
        end else if(en) begin
            t545 <= t544;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t546 <= 0;
        end else if(en) begin
            t546 <= e19;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t547 <= 0;
        end else if(en) begin
            t547 <= f19;
        end
    end
    assign t548 = ($signed(t546) * $signed(t547));
    always @(posedge clock) begin
        if(reset) begin
            t549 <= 0;
        end else if(en) begin
            t549 <= t548;
        end
    end
    assign t550 = ($signed(t549) + $signed(t545));
    always @(posedge clock) begin
        if(reset) begin
            t551 <= 0;
        end else if(en) begin
            t551 <= t550;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t552 <= 0;
        end else if(en) begin
            t552 <= e20;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t553 <= 0;
        end else if(en) begin
            t553 <= f20;
        end
    end
    assign t554 = ($signed(t552) * $signed(t553));
    always @(posedge clock) begin
        if(reset) begin
            t555 <= 0;
        end else if(en) begin
            t555 <= t554;
        end
    end
    assign t556 = ($signed(t555) + $signed(t551));
    always @(posedge clock) begin
        if(reset) begin
            t557 <= 0;
        end else if(en) begin
            t557 <= t556;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t558 <= 0;
        end else if(en) begin
            t558 <= e21;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t559 <= 0;
        end else if(en) begin
            t559 <= f21;
        end
    end
    assign t560 = ($signed(t558) * $signed(t559));
    always @(posedge clock) begin
        if(reset) begin
            t561 <= 0;
        end else if(en) begin
            t561 <= t560;
        end
    end
    assign t562 = ($signed(t561) + $signed(t557));
    always @(posedge clock) begin
        if(reset) begin
            t563 <= 0;
        end else if(en) begin
            t563 <= t562;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t564 <= 0;
        end else if(en) begin
            t564 <= e22;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t565 <= 0;
        end else if(en) begin
            t565 <= f22;
        end
    end
    assign t566 = ($signed(t564) * $signed(t565));
    always @(posedge clock) begin
        if(reset) begin
            t567 <= 0;
        end else if(en) begin
            t567 <= t566;
        end
    end
    assign t568 = ($signed(t567) + $signed(t563));
    always @(posedge clock) begin
        if(reset) begin
            t569 <= 0;
        end else if(en) begin
            t569 <= t568;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t570 <= 0;
        end else if(en) begin
            t570 <= e23;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t571 <= 0;
        end else if(en) begin
            t571 <= f23;
        end
    end
    assign t572 = ($signed(t570) * $signed(t571));
    always @(posedge clock) begin
        if(reset) begin
            t573 <= 0;
        end else if(en) begin
            t573 <= t572;
        end
    end
    assign t574 = ($signed(t573) + $signed(t569));
    always @(posedge clock) begin
        if(reset) begin
            t575 <= 0;
        end else if(en) begin
            t575 <= t574;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t576 <= 0;
        end else if(en) begin
            t576 <= e24;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t577 <= 0;
        end else if(en) begin
            t577 <= f24;
        end
    end
    assign t578 = ($signed(t576) * $signed(t577));
    always @(posedge clock) begin
        if(reset) begin
            t579 <= 0;
        end else if(en) begin
            t579 <= t578;
        end
    end
    assign t580 = ($signed(t579) + $signed(t575));
    always @(posedge clock) begin
        if(reset) begin
            t581 <= 0;
        end else if(en) begin
            t581 <= t580;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t582 <= 0;
        end else if(en) begin
            t582 <= e25;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t583 <= 0;
        end else if(en) begin
            t583 <= f25;
        end
    end
    assign t584 = ($signed(t582) * $signed(t583));
    always @(posedge clock) begin
        if(reset) begin
            t585 <= 0;
        end else if(en) begin
            t585 <= t584;
        end
    end
    assign t586 = ($signed(t585) + $signed(t581));
    always @(posedge clock) begin
        if(reset) begin
            t587 <= 0;
        end else if(en) begin
            t587 <= t586;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t588 <= 0;
        end else if(en) begin
            t588 <= e26;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t589 <= 0;
        end else if(en) begin
            t589 <= f26;
        end
    end
    assign t590 = ($signed(t588) * $signed(t589));
    always @(posedge clock) begin
        if(reset) begin
            t591 <= 0;
        end else if(en) begin
            t591 <= t590;
        end
    end
    assign t592 = ($signed(t591) + $signed(t587));
    always @(posedge clock) begin
        if(reset) begin
            t593 <= 0;
        end else if(en) begin
            t593 <= t592;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t594 <= 0;
        end else if(en) begin
            t594 <= e27;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t595 <= 0;
        end else if(en) begin
            t595 <= f27;
        end
    end
    assign t596 = ($signed(t594) * $signed(t595));
    always @(posedge clock) begin
        if(reset) begin
            t597 <= 0;
        end else if(en) begin
            t597 <= t596;
        end
    end
    assign t598 = ($signed(t597) + $signed(t593));
    always @(posedge clock) begin
        if(reset) begin
            t599 <= 0;
        end else if(en) begin
            t599 <= t598;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t600 <= 0;
        end else if(en) begin
            t600 <= e28;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t601 <= 0;
        end else if(en) begin
            t601 <= f28;
        end
    end
    assign t602 = ($signed(t600) * $signed(t601));
    always @(posedge clock) begin
        if(reset) begin
            t603 <= 0;
        end else if(en) begin
            t603 <= t602;
        end
    end
    assign t604 = ($signed(t603) + $signed(t599));
    always @(posedge clock) begin
        if(reset) begin
            t605 <= 0;
        end else if(en) begin
            t605 <= t604;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t606 <= 0;
        end else if(en) begin
            t606 <= e29;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t607 <= 0;
        end else if(en) begin
            t607 <= f29;
        end
    end
    assign t608 = ($signed(t606) * $signed(t607));
    always @(posedge clock) begin
        if(reset) begin
            t609 <= 0;
        end else if(en) begin
            t609 <= t608;
        end
    end
    assign t610 = ($signed(t609) + $signed(t605));
    always @(posedge clock) begin
        if(reset) begin
            t611 <= 0;
        end else if(en) begin
            t611 <= t610;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t612 <= 0;
        end else if(en) begin
            t612 <= e30;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t613 <= 0;
        end else if(en) begin
            t613 <= f30;
        end
    end
    assign t614 = ($signed(t612) * $signed(t613));
    always @(posedge clock) begin
        if(reset) begin
            t615 <= 0;
        end else if(en) begin
            t615 <= t614;
        end
    end
    assign t616 = ($signed(t615) + $signed(t611));
    always @(posedge clock) begin
        if(reset) begin
            t617 <= 0;
        end else if(en) begin
            t617 <= t616;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t618 <= 0;
        end else if(en) begin
            t618 <= e31;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t619 <= 0;
        end else if(en) begin
            t619 <= f31;
        end
    end
    assign t620 = ($signed(t618) * $signed(t619));
    always @(posedge clock) begin
        if(reset) begin
            t621 <= 0;
        end else if(en) begin
            t621 <= t620;
        end
    end
    assign t622 = ($signed(t621) + $signed(t617));
    always @(posedge clock) begin
        if(reset) begin
            t623 <= 0;
        end else if(en) begin
            t623 <= t622;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t624 <= 0;
        end else if(en) begin
            t624 <= e32;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t625 <= 0;
        end else if(en) begin
            t625 <= f32;
        end
    end
    assign t626 = ($signed(t624) * $signed(t625));
    always @(posedge clock) begin
        if(reset) begin
            t627 <= 0;
        end else if(en) begin
            t627 <= t626;
        end
    end
    assign t628 = ($signed(t627) + $signed(t623));
    always @(posedge clock) begin
        if(reset) begin
            t629 <= 0;
        end else if(en) begin
            t629 <= t628;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t630 <= 0;
        end else if(en) begin
            t630 <= e33;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t631 <= 0;
        end else if(en) begin
            t631 <= f33;
        end
    end
    assign t632 = ($signed(t630) * $signed(t631));
    always @(posedge clock) begin
        if(reset) begin
            t633 <= 0;
        end else if(en) begin
            t633 <= t632;
        end
    end
    assign t634 = ($signed(t633) + $signed(t629));
    always @(posedge clock) begin
        if(reset) begin
            t635 <= 0;
        end else if(en) begin
            t635 <= t634;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t636 <= 0;
        end else if(en) begin
            t636 <= e34;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t637 <= 0;
        end else if(en) begin
            t637 <= f34;
        end
    end
    assign t638 = ($signed(t636) * $signed(t637));
    always @(posedge clock) begin
        if(reset) begin
            t639 <= 0;
        end else if(en) begin
            t639 <= t638;
        end
    end
    assign t640 = ($signed(t639) + $signed(t635));
    always @(posedge clock) begin
        if(reset) begin
            t641 <= 0;
        end else if(en) begin
            t641 <= t640;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t642 <= 0;
        end else if(en) begin
            t642 <= e35;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t643 <= 0;
        end else if(en) begin
            t643 <= f35;
        end
    end
    assign t644 = ($signed(t642) * $signed(t643));
    always @(posedge clock) begin
        if(reset) begin
            t645 <= 0;
        end else if(en) begin
            t645 <= t644;
        end
    end
    assign t646 = ($signed(t645) + $signed(t641));
    always @(posedge clock) begin
        if(reset) begin
            x <= 0;
        end else if(en) begin
            x <= t646;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t648 <= 0;
        end else if(en) begin
            t648 <= g0;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t649 <= 0;
        end else if(en) begin
            t649 <= h0;
        end
    end
    assign t650 = ($signed(t648) * $signed(t649));
    always @(posedge clock) begin
        if(reset) begin
            t651 <= 0;
        end else if(en) begin
            t651 <= t650;
        end
    end
    assign t652 = ($signed(t651) + $signed(p));
    always @(posedge clock) begin
        if(reset) begin
            t653 <= 0;
        end else if(en) begin
            t653 <= t652;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t654 <= 0;
        end else if(en) begin
            t654 <= g1;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t655 <= 0;
        end else if(en) begin
            t655 <= h1;
        end
    end
    assign t656 = ($signed(t654) * $signed(t655));
    always @(posedge clock) begin
        if(reset) begin
            t657 <= 0;
        end else if(en) begin
            t657 <= t656;
        end
    end
    assign t658 = ($signed(t657) + $signed(t653));
    always @(posedge clock) begin
        if(reset) begin
            t659 <= 0;
        end else if(en) begin
            t659 <= t658;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t660 <= 0;
        end else if(en) begin
            t660 <= g2;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t661 <= 0;
        end else if(en) begin
            t661 <= h2;
        end
    end
    assign t662 = ($signed(t660) * $signed(t661));
    always @(posedge clock) begin
        if(reset) begin
            t663 <= 0;
        end else if(en) begin
            t663 <= t662;
        end
    end
    assign t664 = ($signed(t663) + $signed(t659));
    always @(posedge clock) begin
        if(reset) begin
            t665 <= 0;
        end else if(en) begin
            t665 <= t664;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t666 <= 0;
        end else if(en) begin
            t666 <= g3;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t667 <= 0;
        end else if(en) begin
            t667 <= h3;
        end
    end
    assign t668 = ($signed(t666) * $signed(t667));
    always @(posedge clock) begin
        if(reset) begin
            t669 <= 0;
        end else if(en) begin
            t669 <= t668;
        end
    end
    assign t670 = ($signed(t669) + $signed(t665));
    always @(posedge clock) begin
        if(reset) begin
            t671 <= 0;
        end else if(en) begin
            t671 <= t670;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t672 <= 0;
        end else if(en) begin
            t672 <= g4;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t673 <= 0;
        end else if(en) begin
            t673 <= h4;
        end
    end
    assign t674 = ($signed(t672) * $signed(t673));
    always @(posedge clock) begin
        if(reset) begin
            t675 <= 0;
        end else if(en) begin
            t675 <= t674;
        end
    end
    assign t676 = ($signed(t675) + $signed(t671));
    always @(posedge clock) begin
        if(reset) begin
            t677 <= 0;
        end else if(en) begin
            t677 <= t676;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t678 <= 0;
        end else if(en) begin
            t678 <= g5;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t679 <= 0;
        end else if(en) begin
            t679 <= h5;
        end
    end
    assign t680 = ($signed(t678) * $signed(t679));
    always @(posedge clock) begin
        if(reset) begin
            t681 <= 0;
        end else if(en) begin
            t681 <= t680;
        end
    end
    assign t682 = ($signed(t681) + $signed(t677));
    always @(posedge clock) begin
        if(reset) begin
            t683 <= 0;
        end else if(en) begin
            t683 <= t682;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t684 <= 0;
        end else if(en) begin
            t684 <= g6;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t685 <= 0;
        end else if(en) begin
            t685 <= h6;
        end
    end
    assign t686 = ($signed(t684) * $signed(t685));
    always @(posedge clock) begin
        if(reset) begin
            t687 <= 0;
        end else if(en) begin
            t687 <= t686;
        end
    end
    assign t688 = ($signed(t687) + $signed(t683));
    always @(posedge clock) begin
        if(reset) begin
            t689 <= 0;
        end else if(en) begin
            t689 <= t688;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t690 <= 0;
        end else if(en) begin
            t690 <= g7;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t691 <= 0;
        end else if(en) begin
            t691 <= h7;
        end
    end
    assign t692 = ($signed(t690) * $signed(t691));
    always @(posedge clock) begin
        if(reset) begin
            t693 <= 0;
        end else if(en) begin
            t693 <= t692;
        end
    end
    assign t694 = ($signed(t693) + $signed(t689));
    always @(posedge clock) begin
        if(reset) begin
            t695 <= 0;
        end else if(en) begin
            t695 <= t694;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t696 <= 0;
        end else if(en) begin
            t696 <= g8;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t697 <= 0;
        end else if(en) begin
            t697 <= h8;
        end
    end
    assign t698 = ($signed(t696) * $signed(t697));
    always @(posedge clock) begin
        if(reset) begin
            t699 <= 0;
        end else if(en) begin
            t699 <= t698;
        end
    end
    assign t700 = ($signed(t699) + $signed(t695));
    always @(posedge clock) begin
        if(reset) begin
            t701 <= 0;
        end else if(en) begin
            t701 <= t700;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t702 <= 0;
        end else if(en) begin
            t702 <= g9;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t703 <= 0;
        end else if(en) begin
            t703 <= h9;
        end
    end
    assign t704 = ($signed(t702) * $signed(t703));
    always @(posedge clock) begin
        if(reset) begin
            t705 <= 0;
        end else if(en) begin
            t705 <= t704;
        end
    end
    assign t706 = ($signed(t705) + $signed(t701));
    always @(posedge clock) begin
        if(reset) begin
            t707 <= 0;
        end else if(en) begin
            t707 <= t706;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t708 <= 0;
        end else if(en) begin
            t708 <= g10;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t709 <= 0;
        end else if(en) begin
            t709 <= h10;
        end
    end
    assign t710 = ($signed(t708) * $signed(t709));
    always @(posedge clock) begin
        if(reset) begin
            t711 <= 0;
        end else if(en) begin
            t711 <= t710;
        end
    end
    assign t712 = ($signed(t711) + $signed(t707));
    always @(posedge clock) begin
        if(reset) begin
            t713 <= 0;
        end else if(en) begin
            t713 <= t712;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t714 <= 0;
        end else if(en) begin
            t714 <= g11;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t715 <= 0;
        end else if(en) begin
            t715 <= h11;
        end
    end
    assign t716 = ($signed(t714) * $signed(t715));
    always @(posedge clock) begin
        if(reset) begin
            t717 <= 0;
        end else if(en) begin
            t717 <= t716;
        end
    end
    assign t718 = ($signed(t717) + $signed(t713));
    always @(posedge clock) begin
        if(reset) begin
            t719 <= 0;
        end else if(en) begin
            t719 <= t718;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t720 <= 0;
        end else if(en) begin
            t720 <= g12;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t721 <= 0;
        end else if(en) begin
            t721 <= h12;
        end
    end
    assign t722 = ($signed(t720) * $signed(t721));
    always @(posedge clock) begin
        if(reset) begin
            t723 <= 0;
        end else if(en) begin
            t723 <= t722;
        end
    end
    assign t724 = ($signed(t723) + $signed(t719));
    always @(posedge clock) begin
        if(reset) begin
            t725 <= 0;
        end else if(en) begin
            t725 <= t724;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t726 <= 0;
        end else if(en) begin
            t726 <= g13;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t727 <= 0;
        end else if(en) begin
            t727 <= h13;
        end
    end
    assign t728 = ($signed(t726) * $signed(t727));
    always @(posedge clock) begin
        if(reset) begin
            t729 <= 0;
        end else if(en) begin
            t729 <= t728;
        end
    end
    assign t730 = ($signed(t729) + $signed(t725));
    always @(posedge clock) begin
        if(reset) begin
            t731 <= 0;
        end else if(en) begin
            t731 <= t730;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t732 <= 0;
        end else if(en) begin
            t732 <= g14;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t733 <= 0;
        end else if(en) begin
            t733 <= h14;
        end
    end
    assign t734 = ($signed(t732) * $signed(t733));
    always @(posedge clock) begin
        if(reset) begin
            t735 <= 0;
        end else if(en) begin
            t735 <= t734;
        end
    end
    assign t736 = ($signed(t735) + $signed(t731));
    always @(posedge clock) begin
        if(reset) begin
            t737 <= 0;
        end else if(en) begin
            t737 <= t736;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t738 <= 0;
        end else if(en) begin
            t738 <= g15;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t739 <= 0;
        end else if(en) begin
            t739 <= h15;
        end
    end
    assign t740 = ($signed(t738) * $signed(t739));
    always @(posedge clock) begin
        if(reset) begin
            t741 <= 0;
        end else if(en) begin
            t741 <= t740;
        end
    end
    assign t742 = ($signed(t741) + $signed(t737));
    always @(posedge clock) begin
        if(reset) begin
            t743 <= 0;
        end else if(en) begin
            t743 <= t742;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t744 <= 0;
        end else if(en) begin
            t744 <= g16;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t745 <= 0;
        end else if(en) begin
            t745 <= h16;
        end
    end
    assign t746 = ($signed(t744) * $signed(t745));
    always @(posedge clock) begin
        if(reset) begin
            t747 <= 0;
        end else if(en) begin
            t747 <= t746;
        end
    end
    assign t748 = ($signed(t747) + $signed(t743));
    always @(posedge clock) begin
        if(reset) begin
            t749 <= 0;
        end else if(en) begin
            t749 <= t748;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t750 <= 0;
        end else if(en) begin
            t750 <= g17;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t751 <= 0;
        end else if(en) begin
            t751 <= h17;
        end
    end
    assign t752 = ($signed(t750) * $signed(t751));
    always @(posedge clock) begin
        if(reset) begin
            t753 <= 0;
        end else if(en) begin
            t753 <= t752;
        end
    end
    assign t754 = ($signed(t753) + $signed(t749));
    always @(posedge clock) begin
        if(reset) begin
            t755 <= 0;
        end else if(en) begin
            t755 <= t754;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t756 <= 0;
        end else if(en) begin
            t756 <= g18;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t757 <= 0;
        end else if(en) begin
            t757 <= h18;
        end
    end
    assign t758 = ($signed(t756) * $signed(t757));
    always @(posedge clock) begin
        if(reset) begin
            t759 <= 0;
        end else if(en) begin
            t759 <= t758;
        end
    end
    assign t760 = ($signed(t759) + $signed(t755));
    always @(posedge clock) begin
        if(reset) begin
            t761 <= 0;
        end else if(en) begin
            t761 <= t760;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t762 <= 0;
        end else if(en) begin
            t762 <= g19;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t763 <= 0;
        end else if(en) begin
            t763 <= h19;
        end
    end
    assign t764 = ($signed(t762) * $signed(t763));
    always @(posedge clock) begin
        if(reset) begin
            t765 <= 0;
        end else if(en) begin
            t765 <= t764;
        end
    end
    assign t766 = ($signed(t765) + $signed(t761));
    always @(posedge clock) begin
        if(reset) begin
            t767 <= 0;
        end else if(en) begin
            t767 <= t766;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t768 <= 0;
        end else if(en) begin
            t768 <= g20;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t769 <= 0;
        end else if(en) begin
            t769 <= h20;
        end
    end
    assign t770 = ($signed(t768) * $signed(t769));
    always @(posedge clock) begin
        if(reset) begin
            t771 <= 0;
        end else if(en) begin
            t771 <= t770;
        end
    end
    assign t772 = ($signed(t771) + $signed(t767));
    always @(posedge clock) begin
        if(reset) begin
            t773 <= 0;
        end else if(en) begin
            t773 <= t772;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t774 <= 0;
        end else if(en) begin
            t774 <= g21;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t775 <= 0;
        end else if(en) begin
            t775 <= h21;
        end
    end
    assign t776 = ($signed(t774) * $signed(t775));
    always @(posedge clock) begin
        if(reset) begin
            t777 <= 0;
        end else if(en) begin
            t777 <= t776;
        end
    end
    assign t778 = ($signed(t777) + $signed(t773));
    always @(posedge clock) begin
        if(reset) begin
            t779 <= 0;
        end else if(en) begin
            t779 <= t778;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t780 <= 0;
        end else if(en) begin
            t780 <= g22;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t781 <= 0;
        end else if(en) begin
            t781 <= h22;
        end
    end
    assign t782 = ($signed(t780) * $signed(t781));
    always @(posedge clock) begin
        if(reset) begin
            t783 <= 0;
        end else if(en) begin
            t783 <= t782;
        end
    end
    assign t784 = ($signed(t783) + $signed(t779));
    always @(posedge clock) begin
        if(reset) begin
            t785 <= 0;
        end else if(en) begin
            t785 <= t784;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t786 <= 0;
        end else if(en) begin
            t786 <= g23;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t787 <= 0;
        end else if(en) begin
            t787 <= h23;
        end
    end
    assign t788 = ($signed(t786) * $signed(t787));
    always @(posedge clock) begin
        if(reset) begin
            t789 <= 0;
        end else if(en) begin
            t789 <= t788;
        end
    end
    assign t790 = ($signed(t789) + $signed(t785));
    always @(posedge clock) begin
        if(reset) begin
            t791 <= 0;
        end else if(en) begin
            t791 <= t790;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t792 <= 0;
        end else if(en) begin
            t792 <= g24;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t793 <= 0;
        end else if(en) begin
            t793 <= h24;
        end
    end
    assign t794 = ($signed(t792) * $signed(t793));
    always @(posedge clock) begin
        if(reset) begin
            t795 <= 0;
        end else if(en) begin
            t795 <= t794;
        end
    end
    assign t796 = ($signed(t795) + $signed(t791));
    always @(posedge clock) begin
        if(reset) begin
            t797 <= 0;
        end else if(en) begin
            t797 <= t796;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t798 <= 0;
        end else if(en) begin
            t798 <= g25;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t799 <= 0;
        end else if(en) begin
            t799 <= h25;
        end
    end
    assign t800 = ($signed(t798) * $signed(t799));
    always @(posedge clock) begin
        if(reset) begin
            t801 <= 0;
        end else if(en) begin
            t801 <= t800;
        end
    end
    assign t802 = ($signed(t801) + $signed(t797));
    always @(posedge clock) begin
        if(reset) begin
            t803 <= 0;
        end else if(en) begin
            t803 <= t802;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t804 <= 0;
        end else if(en) begin
            t804 <= g26;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t805 <= 0;
        end else if(en) begin
            t805 <= h26;
        end
    end
    assign t806 = ($signed(t804) * $signed(t805));
    always @(posedge clock) begin
        if(reset) begin
            t807 <= 0;
        end else if(en) begin
            t807 <= t806;
        end
    end
    assign t808 = ($signed(t807) + $signed(t803));
    always @(posedge clock) begin
        if(reset) begin
            t809 <= 0;
        end else if(en) begin
            t809 <= t808;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t810 <= 0;
        end else if(en) begin
            t810 <= g27;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t811 <= 0;
        end else if(en) begin
            t811 <= h27;
        end
    end
    assign t812 = ($signed(t810) * $signed(t811));
    always @(posedge clock) begin
        if(reset) begin
            t813 <= 0;
        end else if(en) begin
            t813 <= t812;
        end
    end
    assign t814 = ($signed(t813) + $signed(t809));
    always @(posedge clock) begin
        if(reset) begin
            t815 <= 0;
        end else if(en) begin
            t815 <= t814;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t816 <= 0;
        end else if(en) begin
            t816 <= g28;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t817 <= 0;
        end else if(en) begin
            t817 <= h28;
        end
    end
    assign t818 = ($signed(t816) * $signed(t817));
    always @(posedge clock) begin
        if(reset) begin
            t819 <= 0;
        end else if(en) begin
            t819 <= t818;
        end
    end
    assign t820 = ($signed(t819) + $signed(t815));
    always @(posedge clock) begin
        if(reset) begin
            t821 <= 0;
        end else if(en) begin
            t821 <= t820;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t822 <= 0;
        end else if(en) begin
            t822 <= g29;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t823 <= 0;
        end else if(en) begin
            t823 <= h29;
        end
    end
    assign t824 = ($signed(t822) * $signed(t823));
    always @(posedge clock) begin
        if(reset) begin
            t825 <= 0;
        end else if(en) begin
            t825 <= t824;
        end
    end
    assign t826 = ($signed(t825) + $signed(t821));
    always @(posedge clock) begin
        if(reset) begin
            t827 <= 0;
        end else if(en) begin
            t827 <= t826;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t828 <= 0;
        end else if(en) begin
            t828 <= g30;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t829 <= 0;
        end else if(en) begin
            t829 <= h30;
        end
    end
    assign t830 = ($signed(t828) * $signed(t829));
    always @(posedge clock) begin
        if(reset) begin
            t831 <= 0;
        end else if(en) begin
            t831 <= t830;
        end
    end
    assign t832 = ($signed(t831) + $signed(t827));
    always @(posedge clock) begin
        if(reset) begin
            t833 <= 0;
        end else if(en) begin
            t833 <= t832;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t834 <= 0;
        end else if(en) begin
            t834 <= g31;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t835 <= 0;
        end else if(en) begin
            t835 <= h31;
        end
    end
    assign t836 = ($signed(t834) * $signed(t835));
    always @(posedge clock) begin
        if(reset) begin
            t837 <= 0;
        end else if(en) begin
            t837 <= t836;
        end
    end
    assign t838 = ($signed(t837) + $signed(t833));
    always @(posedge clock) begin
        if(reset) begin
            t839 <= 0;
        end else if(en) begin
            t839 <= t838;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t840 <= 0;
        end else if(en) begin
            t840 <= g32;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t841 <= 0;
        end else if(en) begin
            t841 <= h32;
        end
    end
    assign t842 = ($signed(t840) * $signed(t841));
    always @(posedge clock) begin
        if(reset) begin
            t843 <= 0;
        end else if(en) begin
            t843 <= t842;
        end
    end
    assign t844 = ($signed(t843) + $signed(t839));
    always @(posedge clock) begin
        if(reset) begin
            t845 <= 0;
        end else if(en) begin
            t845 <= t844;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t846 <= 0;
        end else if(en) begin
            t846 <= g33;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t847 <= 0;
        end else if(en) begin
            t847 <= h33;
        end
    end
    assign t848 = ($signed(t846) * $signed(t847));
    always @(posedge clock) begin
        if(reset) begin
            t849 <= 0;
        end else if(en) begin
            t849 <= t848;
        end
    end
    assign t850 = ($signed(t849) + $signed(t845));
    always @(posedge clock) begin
        if(reset) begin
            t851 <= 0;
        end else if(en) begin
            t851 <= t850;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t852 <= 0;
        end else if(en) begin
            t852 <= g34;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t853 <= 0;
        end else if(en) begin
            t853 <= h34;
        end
    end
    assign t854 = ($signed(t852) * $signed(t853));
    always @(posedge clock) begin
        if(reset) begin
            t855 <= 0;
        end else if(en) begin
            t855 <= t854;
        end
    end
    assign t856 = ($signed(t855) + $signed(t851));
    always @(posedge clock) begin
        if(reset) begin
            t857 <= 0;
        end else if(en) begin
            t857 <= t856;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t858 <= 0;
        end else if(en) begin
            t858 <= g35;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t859 <= 0;
        end else if(en) begin
            t859 <= h35;
        end
    end
    assign t860 = ($signed(t858) * $signed(t859));
    always @(posedge clock) begin
        if(reset) begin
            t861 <= 0;
        end else if(en) begin
            t861 <= t860;
        end
    end
    assign t862 = ($signed(t861) + $signed(t857));
    always @(posedge clock) begin
        if(reset) begin
            y <= 0;
        end else if(en) begin
            y <= t862;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t864 <= 0;
        end else if(en) begin
            t864 <= i0;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t865 <= 0;
        end else if(en) begin
            t865 <= j0;
        end
    end
    assign t866 = ($signed(t864) * $signed(t865));
    always @(posedge clock) begin
        if(reset) begin
            t867 <= 0;
        end else if(en) begin
            t867 <= t866;
        end
    end
    assign t868 = ($signed(t867) + $signed(q));
    always @(posedge clock) begin
        if(reset) begin
            t869 <= 0;
        end else if(en) begin
            t869 <= t868;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t870 <= 0;
        end else if(en) begin
            t870 <= i1;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t871 <= 0;
        end else if(en) begin
            t871 <= j1;
        end
    end
    assign t872 = ($signed(t870) * $signed(t871));
    always @(posedge clock) begin
        if(reset) begin
            t873 <= 0;
        end else if(en) begin
            t873 <= t872;
        end
    end
    assign t874 = ($signed(t873) + $signed(t869));
    always @(posedge clock) begin
        if(reset) begin
            t875 <= 0;
        end else if(en) begin
            t875 <= t874;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t876 <= 0;
        end else if(en) begin
            t876 <= i2;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t877 <= 0;
        end else if(en) begin
            t877 <= j2;
        end
    end
    assign t878 = ($signed(t876) * $signed(t877));
    always @(posedge clock) begin
        if(reset) begin
            t879 <= 0;
        end else if(en) begin
            t879 <= t878;
        end
    end
    assign t880 = ($signed(t879) + $signed(t875));
    always @(posedge clock) begin
        if(reset) begin
            t881 <= 0;
        end else if(en) begin
            t881 <= t880;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t882 <= 0;
        end else if(en) begin
            t882 <= i3;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t883 <= 0;
        end else if(en) begin
            t883 <= j3;
        end
    end
    assign t884 = ($signed(t882) * $signed(t883));
    always @(posedge clock) begin
        if(reset) begin
            t885 <= 0;
        end else if(en) begin
            t885 <= t884;
        end
    end
    assign t886 = ($signed(t885) + $signed(t881));
    always @(posedge clock) begin
        if(reset) begin
            t887 <= 0;
        end else if(en) begin
            t887 <= t886;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t888 <= 0;
        end else if(en) begin
            t888 <= i4;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t889 <= 0;
        end else if(en) begin
            t889 <= j4;
        end
    end
    assign t890 = ($signed(t888) * $signed(t889));
    always @(posedge clock) begin
        if(reset) begin
            t891 <= 0;
        end else if(en) begin
            t891 <= t890;
        end
    end
    assign t892 = ($signed(t891) + $signed(t887));
    always @(posedge clock) begin
        if(reset) begin
            t893 <= 0;
        end else if(en) begin
            t893 <= t892;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t894 <= 0;
        end else if(en) begin
            t894 <= i5;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t895 <= 0;
        end else if(en) begin
            t895 <= j5;
        end
    end
    assign t896 = ($signed(t894) * $signed(t895));
    always @(posedge clock) begin
        if(reset) begin
            t897 <= 0;
        end else if(en) begin
            t897 <= t896;
        end
    end
    assign t898 = ($signed(t897) + $signed(t893));
    always @(posedge clock) begin
        if(reset) begin
            t899 <= 0;
        end else if(en) begin
            t899 <= t898;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t900 <= 0;
        end else if(en) begin
            t900 <= i6;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t901 <= 0;
        end else if(en) begin
            t901 <= j6;
        end
    end
    assign t902 = ($signed(t900) * $signed(t901));
    always @(posedge clock) begin
        if(reset) begin
            t903 <= 0;
        end else if(en) begin
            t903 <= t902;
        end
    end
    assign t904 = ($signed(t903) + $signed(t899));
    always @(posedge clock) begin
        if(reset) begin
            t905 <= 0;
        end else if(en) begin
            t905 <= t904;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t906 <= 0;
        end else if(en) begin
            t906 <= i7;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t907 <= 0;
        end else if(en) begin
            t907 <= j7;
        end
    end
    assign t908 = ($signed(t906) * $signed(t907));
    always @(posedge clock) begin
        if(reset) begin
            t909 <= 0;
        end else if(en) begin
            t909 <= t908;
        end
    end
    assign t910 = ($signed(t909) + $signed(t905));
    always @(posedge clock) begin
        if(reset) begin
            t911 <= 0;
        end else if(en) begin
            t911 <= t910;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t912 <= 0;
        end else if(en) begin
            t912 <= i8;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t913 <= 0;
        end else if(en) begin
            t913 <= j8;
        end
    end
    assign t914 = ($signed(t912) * $signed(t913));
    always @(posedge clock) begin
        if(reset) begin
            t915 <= 0;
        end else if(en) begin
            t915 <= t914;
        end
    end
    assign t916 = ($signed(t915) + $signed(t911));
    always @(posedge clock) begin
        if(reset) begin
            t917 <= 0;
        end else if(en) begin
            t917 <= t916;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t918 <= 0;
        end else if(en) begin
            t918 <= i9;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t919 <= 0;
        end else if(en) begin
            t919 <= j9;
        end
    end
    assign t920 = ($signed(t918) * $signed(t919));
    always @(posedge clock) begin
        if(reset) begin
            t921 <= 0;
        end else if(en) begin
            t921 <= t920;
        end
    end
    assign t922 = ($signed(t921) + $signed(t917));
    always @(posedge clock) begin
        if(reset) begin
            t923 <= 0;
        end else if(en) begin
            t923 <= t922;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t924 <= 0;
        end else if(en) begin
            t924 <= i10;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t925 <= 0;
        end else if(en) begin
            t925 <= j10;
        end
    end
    assign t926 = ($signed(t924) * $signed(t925));
    always @(posedge clock) begin
        if(reset) begin
            t927 <= 0;
        end else if(en) begin
            t927 <= t926;
        end
    end
    assign t928 = ($signed(t927) + $signed(t923));
    always @(posedge clock) begin
        if(reset) begin
            t929 <= 0;
        end else if(en) begin
            t929 <= t928;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t930 <= 0;
        end else if(en) begin
            t930 <= i11;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t931 <= 0;
        end else if(en) begin
            t931 <= j11;
        end
    end
    assign t932 = ($signed(t930) * $signed(t931));
    always @(posedge clock) begin
        if(reset) begin
            t933 <= 0;
        end else if(en) begin
            t933 <= t932;
        end
    end
    assign t934 = ($signed(t933) + $signed(t929));
    always @(posedge clock) begin
        if(reset) begin
            t935 <= 0;
        end else if(en) begin
            t935 <= t934;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t936 <= 0;
        end else if(en) begin
            t936 <= i12;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t937 <= 0;
        end else if(en) begin
            t937 <= j12;
        end
    end
    assign t938 = ($signed(t936) * $signed(t937));
    always @(posedge clock) begin
        if(reset) begin
            t939 <= 0;
        end else if(en) begin
            t939 <= t938;
        end
    end
    assign t940 = ($signed(t939) + $signed(t935));
    always @(posedge clock) begin
        if(reset) begin
            t941 <= 0;
        end else if(en) begin
            t941 <= t940;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t942 <= 0;
        end else if(en) begin
            t942 <= i13;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t943 <= 0;
        end else if(en) begin
            t943 <= j13;
        end
    end
    assign t944 = ($signed(t942) * $signed(t943));
    always @(posedge clock) begin
        if(reset) begin
            t945 <= 0;
        end else if(en) begin
            t945 <= t944;
        end
    end
    assign t946 = ($signed(t945) + $signed(t941));
    always @(posedge clock) begin
        if(reset) begin
            t947 <= 0;
        end else if(en) begin
            t947 <= t946;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t948 <= 0;
        end else if(en) begin
            t948 <= i14;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t949 <= 0;
        end else if(en) begin
            t949 <= j14;
        end
    end
    assign t950 = ($signed(t948) * $signed(t949));
    always @(posedge clock) begin
        if(reset) begin
            t951 <= 0;
        end else if(en) begin
            t951 <= t950;
        end
    end
    assign t952 = ($signed(t951) + $signed(t947));
    always @(posedge clock) begin
        if(reset) begin
            t953 <= 0;
        end else if(en) begin
            t953 <= t952;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t954 <= 0;
        end else if(en) begin
            t954 <= i15;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t955 <= 0;
        end else if(en) begin
            t955 <= j15;
        end
    end
    assign t956 = ($signed(t954) * $signed(t955));
    always @(posedge clock) begin
        if(reset) begin
            t957 <= 0;
        end else if(en) begin
            t957 <= t956;
        end
    end
    assign t958 = ($signed(t957) + $signed(t953));
    always @(posedge clock) begin
        if(reset) begin
            t959 <= 0;
        end else if(en) begin
            t959 <= t958;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t960 <= 0;
        end else if(en) begin
            t960 <= i16;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t961 <= 0;
        end else if(en) begin
            t961 <= j16;
        end
    end
    assign t962 = ($signed(t960) * $signed(t961));
    always @(posedge clock) begin
        if(reset) begin
            t963 <= 0;
        end else if(en) begin
            t963 <= t962;
        end
    end
    assign t964 = ($signed(t963) + $signed(t959));
    always @(posedge clock) begin
        if(reset) begin
            t965 <= 0;
        end else if(en) begin
            t965 <= t964;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t966 <= 0;
        end else if(en) begin
            t966 <= i17;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t967 <= 0;
        end else if(en) begin
            t967 <= j17;
        end
    end
    assign t968 = ($signed(t966) * $signed(t967));
    always @(posedge clock) begin
        if(reset) begin
            t969 <= 0;
        end else if(en) begin
            t969 <= t968;
        end
    end
    assign t970 = ($signed(t969) + $signed(t965));
    always @(posedge clock) begin
        if(reset) begin
            t971 <= 0;
        end else if(en) begin
            t971 <= t970;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t972 <= 0;
        end else if(en) begin
            t972 <= i18;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t973 <= 0;
        end else if(en) begin
            t973 <= j18;
        end
    end
    assign t974 = ($signed(t972) * $signed(t973));
    always @(posedge clock) begin
        if(reset) begin
            t975 <= 0;
        end else if(en) begin
            t975 <= t974;
        end
    end
    assign t976 = ($signed(t975) + $signed(t971));
    always @(posedge clock) begin
        if(reset) begin
            t977 <= 0;
        end else if(en) begin
            t977 <= t976;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t978 <= 0;
        end else if(en) begin
            t978 <= i19;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t979 <= 0;
        end else if(en) begin
            t979 <= j19;
        end
    end
    assign t980 = ($signed(t978) * $signed(t979));
    always @(posedge clock) begin
        if(reset) begin
            t981 <= 0;
        end else if(en) begin
            t981 <= t980;
        end
    end
    assign t982 = ($signed(t981) + $signed(t977));
    always @(posedge clock) begin
        if(reset) begin
            t983 <= 0;
        end else if(en) begin
            t983 <= t982;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t984 <= 0;
        end else if(en) begin
            t984 <= i20;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t985 <= 0;
        end else if(en) begin
            t985 <= j20;
        end
    end
    assign t986 = ($signed(t984) * $signed(t985));
    always @(posedge clock) begin
        if(reset) begin
            t987 <= 0;
        end else if(en) begin
            t987 <= t986;
        end
    end
    assign t988 = ($signed(t987) + $signed(t983));
    always @(posedge clock) begin
        if(reset) begin
            t989 <= 0;
        end else if(en) begin
            t989 <= t988;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t990 <= 0;
        end else if(en) begin
            t990 <= i21;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t991 <= 0;
        end else if(en) begin
            t991 <= j21;
        end
    end
    assign t992 = ($signed(t990) * $signed(t991));
    always @(posedge clock) begin
        if(reset) begin
            t993 <= 0;
        end else if(en) begin
            t993 <= t992;
        end
    end
    assign t994 = ($signed(t993) + $signed(t989));
    always @(posedge clock) begin
        if(reset) begin
            t995 <= 0;
        end else if(en) begin
            t995 <= t994;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t996 <= 0;
        end else if(en) begin
            t996 <= i22;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t997 <= 0;
        end else if(en) begin
            t997 <= j22;
        end
    end
    assign t998 = ($signed(t996) * $signed(t997));
    always @(posedge clock) begin
        if(reset) begin
            t999 <= 0;
        end else if(en) begin
            t999 <= t998;
        end
    end
    assign t1000 = ($signed(t999) + $signed(t995));
    always @(posedge clock) begin
        if(reset) begin
            t1001 <= 0;
        end else if(en) begin
            t1001 <= t1000;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t1002 <= 0;
        end else if(en) begin
            t1002 <= i23;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t1003 <= 0;
        end else if(en) begin
            t1003 <= j23;
        end
    end
    assign t1004 = ($signed(t1002) * $signed(t1003));
    always @(posedge clock) begin
        if(reset) begin
            t1005 <= 0;
        end else if(en) begin
            t1005 <= t1004;
        end
    end
    assign t1006 = ($signed(t1005) + $signed(t1001));
    always @(posedge clock) begin
        if(reset) begin
            t1007 <= 0;
        end else if(en) begin
            t1007 <= t1006;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t1008 <= 0;
        end else if(en) begin
            t1008 <= i24;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t1009 <= 0;
        end else if(en) begin
            t1009 <= j24;
        end
    end
    assign t1010 = ($signed(t1008) * $signed(t1009));
    always @(posedge clock) begin
        if(reset) begin
            t1011 <= 0;
        end else if(en) begin
            t1011 <= t1010;
        end
    end
    assign t1012 = ($signed(t1011) + $signed(t1007));
    always @(posedge clock) begin
        if(reset) begin
            t1013 <= 0;
        end else if(en) begin
            t1013 <= t1012;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t1014 <= 0;
        end else if(en) begin
            t1014 <= i25;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t1015 <= 0;
        end else if(en) begin
            t1015 <= j25;
        end
    end
    assign t1016 = ($signed(t1014) * $signed(t1015));
    always @(posedge clock) begin
        if(reset) begin
            t1017 <= 0;
        end else if(en) begin
            t1017 <= t1016;
        end
    end
    assign t1018 = ($signed(t1017) + $signed(t1013));
    always @(posedge clock) begin
        if(reset) begin
            t1019 <= 0;
        end else if(en) begin
            t1019 <= t1018;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t1020 <= 0;
        end else if(en) begin
            t1020 <= i26;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t1021 <= 0;
        end else if(en) begin
            t1021 <= j26;
        end
    end
    assign t1022 = ($signed(t1020) * $signed(t1021));
    always @(posedge clock) begin
        if(reset) begin
            t1023 <= 0;
        end else if(en) begin
            t1023 <= t1022;
        end
    end
    assign t1024 = ($signed(t1023) + $signed(t1019));
    always @(posedge clock) begin
        if(reset) begin
            t1025 <= 0;
        end else if(en) begin
            t1025 <= t1024;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t1026 <= 0;
        end else if(en) begin
            t1026 <= i27;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t1027 <= 0;
        end else if(en) begin
            t1027 <= j27;
        end
    end
    assign t1028 = ($signed(t1026) * $signed(t1027));
    always @(posedge clock) begin
        if(reset) begin
            t1029 <= 0;
        end else if(en) begin
            t1029 <= t1028;
        end
    end
    assign t1030 = ($signed(t1029) + $signed(t1025));
    always @(posedge clock) begin
        if(reset) begin
            t1031 <= 0;
        end else if(en) begin
            t1031 <= t1030;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t1032 <= 0;
        end else if(en) begin
            t1032 <= i28;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t1033 <= 0;
        end else if(en) begin
            t1033 <= j28;
        end
    end
    assign t1034 = ($signed(t1032) * $signed(t1033));
    always @(posedge clock) begin
        if(reset) begin
            t1035 <= 0;
        end else if(en) begin
            t1035 <= t1034;
        end
    end
    assign t1036 = ($signed(t1035) + $signed(t1031));
    always @(posedge clock) begin
        if(reset) begin
            t1037 <= 0;
        end else if(en) begin
            t1037 <= t1036;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t1038 <= 0;
        end else if(en) begin
            t1038 <= i29;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t1039 <= 0;
        end else if(en) begin
            t1039 <= j29;
        end
    end
    assign t1040 = ($signed(t1038) * $signed(t1039));
    always @(posedge clock) begin
        if(reset) begin
            t1041 <= 0;
        end else if(en) begin
            t1041 <= t1040;
        end
    end
    assign t1042 = ($signed(t1041) + $signed(t1037));
    always @(posedge clock) begin
        if(reset) begin
            t1043 <= 0;
        end else if(en) begin
            t1043 <= t1042;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t1044 <= 0;
        end else if(en) begin
            t1044 <= i30;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t1045 <= 0;
        end else if(en) begin
            t1045 <= j30;
        end
    end
    assign t1046 = ($signed(t1044) * $signed(t1045));
    always @(posedge clock) begin
        if(reset) begin
            t1047 <= 0;
        end else if(en) begin
            t1047 <= t1046;
        end
    end
    assign t1048 = ($signed(t1047) + $signed(t1043));
    always @(posedge clock) begin
        if(reset) begin
            t1049 <= 0;
        end else if(en) begin
            t1049 <= t1048;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t1050 <= 0;
        end else if(en) begin
            t1050 <= i31;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t1051 <= 0;
        end else if(en) begin
            t1051 <= j31;
        end
    end
    assign t1052 = ($signed(t1050) * $signed(t1051));
    always @(posedge clock) begin
        if(reset) begin
            t1053 <= 0;
        end else if(en) begin
            t1053 <= t1052;
        end
    end
    assign t1054 = ($signed(t1053) + $signed(t1049));
    always @(posedge clock) begin
        if(reset) begin
            t1055 <= 0;
        end else if(en) begin
            t1055 <= t1054;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t1056 <= 0;
        end else if(en) begin
            t1056 <= i32;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t1057 <= 0;
        end else if(en) begin
            t1057 <= j32;
        end
    end
    assign t1058 = ($signed(t1056) * $signed(t1057));
    always @(posedge clock) begin
        if(reset) begin
            t1059 <= 0;
        end else if(en) begin
            t1059 <= t1058;
        end
    end
    assign t1060 = ($signed(t1059) + $signed(t1055));
    always @(posedge clock) begin
        if(reset) begin
            t1061 <= 0;
        end else if(en) begin
            t1061 <= t1060;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t1062 <= 0;
        end else if(en) begin
            t1062 <= i33;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t1063 <= 0;
        end else if(en) begin
            t1063 <= j33;
        end
    end
    assign t1064 = ($signed(t1062) * $signed(t1063));
    always @(posedge clock) begin
        if(reset) begin
            t1065 <= 0;
        end else if(en) begin
            t1065 <= t1064;
        end
    end
    assign t1066 = ($signed(t1065) + $signed(t1061));
    always @(posedge clock) begin
        if(reset) begin
            t1067 <= 0;
        end else if(en) begin
            t1067 <= t1066;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t1068 <= 0;
        end else if(en) begin
            t1068 <= i34;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t1069 <= 0;
        end else if(en) begin
            t1069 <= j34;
        end
    end
    assign t1070 = ($signed(t1068) * $signed(t1069));
    always @(posedge clock) begin
        if(reset) begin
            t1071 <= 0;
        end else if(en) begin
            t1071 <= t1070;
        end
    end
    assign t1072 = ($signed(t1071) + $signed(t1067));
    always @(posedge clock) begin
        if(reset) begin
            t1073 <= 0;
        end else if(en) begin
            t1073 <= t1072;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t1074 <= 0;
        end else if(en) begin
            t1074 <= i35;
        end
    end
    always @(posedge clock) begin
        if(reset) begin
            t1075 <= 0;
        end else if(en) begin
            t1075 <= j35;
        end
    end
    assign t1076 = ($signed(t1074) * $signed(t1075));
    always @(posedge clock) begin
        if(reset) begin
            t1077 <= 0;
        end else if(en) begin
            t1077 <= t1076;
        end
    end
    assign t1078 = ($signed(t1077) + $signed(t1073));
    always @(posedge clock) begin
        if(reset) begin
            z <= 0;
        end else if(en) begin
            z <= t1078;
        end
    end
endmodule
